library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- library SYSTEM_TYPES;
use work.SYSTEM_TYPES.ALL;

-- library CUSTOM_TYPES;
use work.CUSTOM_TYPES.ALL;

-- User defined packages here
-- #### USER-DATA-IMPORTS-START
-- #### USER-DATA-IMPORTS-END

entity sme_intro_export is
    port(
        -- Top-level bus nfa_dfa_Control signals
        nfa_dfa_Control_Valid: out STD_LOGIC;
        nfa_dfa_Control_Reset: out STD_LOGIC;
        nfa_dfa_Control_Length: out STD_LOGIC_VECTOR(31 downto 0);
        nfa_dfa_Control_Array0: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array1: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array2: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array3: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array4: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array5: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array6: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array7: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array8: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array9: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array10: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array11: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array12: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array13: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array14: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array15: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array16: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array17: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array18: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array19: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array20: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array21: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array22: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array23: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array24: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array25: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array26: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array27: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array28: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array29: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array30: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array31: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array32: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array33: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array34: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array35: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array36: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array37: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array38: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array39: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array40: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array41: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array42: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array43: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array44: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array45: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array46: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array47: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array48: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array49: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array50: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array51: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array52: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array53: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array54: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array55: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array56: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array57: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array58: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array59: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array60: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array61: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array62: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array63: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array64: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array65: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array66: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array67: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array68: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array69: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array70: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array71: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array72: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array73: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array74: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array75: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array76: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array77: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array78: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array79: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array80: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array81: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array82: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array83: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array84: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array85: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array86: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array87: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array88: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array89: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array90: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array91: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array92: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array93: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array94: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array95: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array96: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array97: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array98: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array99: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array100: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array101: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array102: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array103: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array104: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array105: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array106: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array107: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array108: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array109: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array110: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array111: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array112: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array113: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array114: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array115: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array116: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array117: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array118: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array119: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array120: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array121: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array122: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array123: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array124: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array125: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array126: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array127: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array128: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array129: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array130: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array131: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array132: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array133: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array134: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array135: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array136: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array137: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array138: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array139: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array140: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array141: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array142: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array143: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array144: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array145: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array146: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array147: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array148: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array149: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array150: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array151: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array152: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array153: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array154: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array155: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array156: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array157: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array158: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array159: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array160: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array161: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array162: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array163: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array164: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array165: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array166: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array167: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array168: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array169: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array170: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array171: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array172: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array173: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array174: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array175: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array176: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array177: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array178: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array179: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array180: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array181: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array182: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array183: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array184: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array185: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array186: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array187: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array188: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array189: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array190: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array191: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array192: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array193: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array194: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array195: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array196: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array197: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array198: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array199: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array200: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array201: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array202: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array203: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array204: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array205: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array206: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array207: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array208: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array209: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array210: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array211: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array212: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array213: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array214: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array215: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array216: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array217: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array218: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array219: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array220: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array221: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array222: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array223: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array224: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array225: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array226: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array227: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array228: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array229: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array230: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array231: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array232: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array233: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array234: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array235: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array236: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array237: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array238: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array239: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array240: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array241: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array242: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array243: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array244: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array245: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array246: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array247: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array248: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array249: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array250: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array251: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array252: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array253: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array254: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array255: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array256: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array257: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array258: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array259: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array260: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array261: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array262: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array263: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array264: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array265: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array266: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array267: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array268: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array269: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array270: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array271: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array272: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array273: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array274: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array275: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array276: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array277: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array278: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array279: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array280: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array281: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array282: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array283: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array284: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array285: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array286: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array287: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array288: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array289: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array290: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array291: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array292: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array293: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array294: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array295: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array296: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array297: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array298: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array299: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array300: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array301: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array302: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array303: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array304: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array305: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array306: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array307: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array308: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array309: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array310: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array311: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array312: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array313: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array314: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array315: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array316: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array317: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array318: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array319: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array320: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array321: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array322: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array323: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array324: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array325: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array326: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array327: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array328: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array329: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array330: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array331: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array332: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array333: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array334: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array335: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array336: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array337: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array338: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array339: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array340: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array341: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array342: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array343: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array344: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array345: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array346: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array347: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array348: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array349: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array350: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array351: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array352: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array353: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array354: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array355: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array356: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array357: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array358: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array359: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array360: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array361: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array362: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array363: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array364: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array365: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array366: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array367: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array368: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array369: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array370: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array371: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array372: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array373: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array374: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array375: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array376: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array377: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array378: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array379: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array380: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array381: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array382: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array383: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array384: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array385: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array386: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array387: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array388: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array389: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array390: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array391: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array392: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array393: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array394: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array395: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array396: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array397: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array398: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array399: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array400: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array401: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array402: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array403: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array404: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array405: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array406: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array407: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array408: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array409: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array410: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array411: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array412: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array413: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array414: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array415: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array416: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array417: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array418: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array419: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array420: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array421: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array422: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array423: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array424: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array425: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array426: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array427: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array428: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array429: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array430: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array431: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array432: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array433: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array434: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array435: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array436: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array437: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array438: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array439: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array440: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array441: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array442: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array443: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array444: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array445: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array446: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array447: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array448: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array449: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array450: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array451: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array452: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array453: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array454: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array455: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array456: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array457: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array458: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array459: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array460: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array461: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array462: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array463: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array464: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array465: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array466: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array467: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array468: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array469: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array470: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array471: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array472: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array473: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array474: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array475: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array476: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array477: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array478: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array479: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array480: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array481: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array482: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array483: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array484: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array485: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array486: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array487: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array488: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array489: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array490: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array491: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array492: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array493: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array494: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array495: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array496: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array497: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array498: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array499: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array500: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array501: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array502: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array503: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array504: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array505: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array506: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array507: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array508: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array509: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array510: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array511: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array512: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array513: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array514: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array515: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array516: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array517: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array518: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array519: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array520: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array521: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array522: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array523: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array524: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array525: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array526: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array527: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array528: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array529: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array530: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array531: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array532: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array533: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array534: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array535: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array536: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array537: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array538: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array539: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array540: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array541: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array542: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array543: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array544: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array545: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array546: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array547: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array548: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array549: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array550: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array551: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array552: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array553: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array554: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array555: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array556: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array557: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array558: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array559: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array560: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array561: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array562: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array563: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array564: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array565: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array566: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array567: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array568: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array569: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array570: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array571: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array572: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array573: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array574: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array575: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array576: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array577: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array578: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array579: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array580: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array581: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array582: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array583: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array584: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array585: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array586: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array587: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array588: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array589: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array590: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array591: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array592: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array593: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array594: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array595: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array596: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array597: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array598: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array599: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array600: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array601: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array602: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array603: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array604: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array605: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array606: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array607: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array608: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array609: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array610: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array611: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array612: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array613: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array614: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array615: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array616: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array617: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array618: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array619: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array620: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array621: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array622: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array623: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array624: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array625: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array626: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array627: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array628: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array629: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array630: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array631: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array632: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array633: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array634: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array635: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array636: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array637: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array638: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array639: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array640: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array641: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array642: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array643: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array644: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array645: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array646: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array647: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array648: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array649: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array650: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array651: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array652: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array653: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array654: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array655: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array656: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array657: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array658: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array659: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array660: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array661: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array662: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array663: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array664: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array665: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array666: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array667: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array668: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array669: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array670: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array671: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array672: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array673: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array674: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array675: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array676: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array677: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array678: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array679: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array680: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array681: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array682: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array683: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array684: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array685: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array686: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array687: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array688: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array689: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array690: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array691: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array692: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array693: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array694: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array695: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array696: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array697: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array698: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array699: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array700: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array701: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array702: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array703: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array704: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array705: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array706: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array707: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array708: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array709: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array710: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array711: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array712: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array713: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array714: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array715: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array716: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array717: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array718: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array719: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array720: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array721: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array722: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array723: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array724: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array725: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array726: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array727: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array728: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array729: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array730: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array731: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array732: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array733: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array734: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array735: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array736: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array737: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array738: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array739: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array740: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array741: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array742: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array743: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array744: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array745: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array746: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array747: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array748: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array749: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array750: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array751: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array752: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array753: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array754: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array755: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array756: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array757: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array758: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array759: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array760: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array761: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array762: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array763: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array764: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array765: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array766: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array767: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array768: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array769: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array770: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array771: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array772: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array773: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array774: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array775: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array776: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array777: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array778: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array779: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array780: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array781: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array782: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array783: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array784: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array785: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array786: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array787: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array788: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array789: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array790: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array791: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array792: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array793: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array794: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array795: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array796: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array797: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array798: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array799: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array800: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array801: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array802: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array803: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array804: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array805: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array806: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array807: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array808: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array809: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array810: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array811: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array812: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array813: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array814: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array815: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array816: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array817: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array818: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array819: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array820: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array821: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array822: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array823: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array824: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array825: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array826: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array827: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array828: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array829: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array830: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array831: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array832: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array833: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array834: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array835: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array836: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array837: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array838: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array839: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array840: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array841: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array842: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array843: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array844: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array845: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array846: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array847: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array848: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array849: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array850: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array851: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array852: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array853: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array854: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array855: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array856: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array857: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array858: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array859: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array860: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array861: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array862: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array863: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array864: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array865: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array866: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array867: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array868: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array869: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array870: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array871: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array872: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array873: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array874: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array875: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array876: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array877: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array878: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array879: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array880: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array881: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array882: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array883: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array884: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array885: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array886: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array887: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array888: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array889: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array890: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array891: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array892: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array893: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array894: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array895: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array896: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array897: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array898: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array899: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array900: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array901: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array902: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array903: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array904: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array905: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array906: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array907: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array908: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array909: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array910: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array911: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array912: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array913: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array914: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array915: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array916: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array917: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array918: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array919: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array920: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array921: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array922: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array923: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array924: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array925: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array926: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array927: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array928: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array929: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array930: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array931: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array932: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array933: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array934: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array935: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array936: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array937: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array938: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array939: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array940: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array941: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array942: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array943: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array944: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array945: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array946: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array947: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array948: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array949: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array950: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array951: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array952: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array953: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array954: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array955: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array956: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array957: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array958: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array959: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array960: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array961: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array962: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array963: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array964: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array965: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array966: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array967: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array968: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array969: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array970: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array971: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array972: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array973: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array974: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array975: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array976: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array977: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array978: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array979: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array980: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array981: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array982: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array983: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array984: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array985: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array986: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array987: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array988: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array989: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array990: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array991: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array992: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array993: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array994: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array995: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array996: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array997: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array998: out STD_LOGIC_VECTOR(7 downto 0);
        nfa_dfa_Control_Array999: out STD_LOGIC_VECTOR(7 downto 0);

        -- Top-level bus nfa_dfa_Traversal signals
        nfa_dfa_Traversal_Valid: in STD_LOGIC;

        -- User defined signals here
        -- #### USER-DATA-ENTITYSIGNALS-START
        -- #### USER-DATA-ENTITYSIGNALS-END

        -- Enable signal
        ENB : in STD_LOGIC;

        -- Reset signal
        RST : in STD_LOGIC;

        -- Finished signal
        FIN : out Std_logic;

        -- Clock signal
        CLK : in STD_LOGIC
    );
end sme_intro_export;

architecture RTL of sme_intro_export is

    -- User defined signals here
    -- #### USER-DATA-SIGNALS-START
    -- #### USER-DATA-SIGNALS-END

    -- Intermediate conversion signal to convert internal types to external ones
    signal tmp_nfa_dfa_Control_Length : T_SYSTEM_INT32;
    signal tmp_nfa_dfa_Control_Array : nfa_dfa_Control_Array_type;

begin

    -- Carry converted signals from entity to wrapped outputs
    nfa_dfa_Control_Length <= std_logic_vector(tmp_nfa_dfa_Control_Length);
    nfa_dfa_Control_Array0 <= std_logic_vector(tmp_nfa_dfa_Control_Array(0));
    nfa_dfa_Control_Array1 <= std_logic_vector(tmp_nfa_dfa_Control_Array(1));
    nfa_dfa_Control_Array2 <= std_logic_vector(tmp_nfa_dfa_Control_Array(2));
    nfa_dfa_Control_Array3 <= std_logic_vector(tmp_nfa_dfa_Control_Array(3));
    nfa_dfa_Control_Array4 <= std_logic_vector(tmp_nfa_dfa_Control_Array(4));
    nfa_dfa_Control_Array5 <= std_logic_vector(tmp_nfa_dfa_Control_Array(5));
    nfa_dfa_Control_Array6 <= std_logic_vector(tmp_nfa_dfa_Control_Array(6));
    nfa_dfa_Control_Array7 <= std_logic_vector(tmp_nfa_dfa_Control_Array(7));
    nfa_dfa_Control_Array8 <= std_logic_vector(tmp_nfa_dfa_Control_Array(8));
    nfa_dfa_Control_Array9 <= std_logic_vector(tmp_nfa_dfa_Control_Array(9));
    nfa_dfa_Control_Array10 <= std_logic_vector(tmp_nfa_dfa_Control_Array(10));
    nfa_dfa_Control_Array11 <= std_logic_vector(tmp_nfa_dfa_Control_Array(11));
    nfa_dfa_Control_Array12 <= std_logic_vector(tmp_nfa_dfa_Control_Array(12));
    nfa_dfa_Control_Array13 <= std_logic_vector(tmp_nfa_dfa_Control_Array(13));
    nfa_dfa_Control_Array14 <= std_logic_vector(tmp_nfa_dfa_Control_Array(14));
    nfa_dfa_Control_Array15 <= std_logic_vector(tmp_nfa_dfa_Control_Array(15));
    nfa_dfa_Control_Array16 <= std_logic_vector(tmp_nfa_dfa_Control_Array(16));
    nfa_dfa_Control_Array17 <= std_logic_vector(tmp_nfa_dfa_Control_Array(17));
    nfa_dfa_Control_Array18 <= std_logic_vector(tmp_nfa_dfa_Control_Array(18));
    nfa_dfa_Control_Array19 <= std_logic_vector(tmp_nfa_dfa_Control_Array(19));
    nfa_dfa_Control_Array20 <= std_logic_vector(tmp_nfa_dfa_Control_Array(20));
    nfa_dfa_Control_Array21 <= std_logic_vector(tmp_nfa_dfa_Control_Array(21));
    nfa_dfa_Control_Array22 <= std_logic_vector(tmp_nfa_dfa_Control_Array(22));
    nfa_dfa_Control_Array23 <= std_logic_vector(tmp_nfa_dfa_Control_Array(23));
    nfa_dfa_Control_Array24 <= std_logic_vector(tmp_nfa_dfa_Control_Array(24));
    nfa_dfa_Control_Array25 <= std_logic_vector(tmp_nfa_dfa_Control_Array(25));
    nfa_dfa_Control_Array26 <= std_logic_vector(tmp_nfa_dfa_Control_Array(26));
    nfa_dfa_Control_Array27 <= std_logic_vector(tmp_nfa_dfa_Control_Array(27));
    nfa_dfa_Control_Array28 <= std_logic_vector(tmp_nfa_dfa_Control_Array(28));
    nfa_dfa_Control_Array29 <= std_logic_vector(tmp_nfa_dfa_Control_Array(29));
    nfa_dfa_Control_Array30 <= std_logic_vector(tmp_nfa_dfa_Control_Array(30));
    nfa_dfa_Control_Array31 <= std_logic_vector(tmp_nfa_dfa_Control_Array(31));
    nfa_dfa_Control_Array32 <= std_logic_vector(tmp_nfa_dfa_Control_Array(32));
    nfa_dfa_Control_Array33 <= std_logic_vector(tmp_nfa_dfa_Control_Array(33));
    nfa_dfa_Control_Array34 <= std_logic_vector(tmp_nfa_dfa_Control_Array(34));
    nfa_dfa_Control_Array35 <= std_logic_vector(tmp_nfa_dfa_Control_Array(35));
    nfa_dfa_Control_Array36 <= std_logic_vector(tmp_nfa_dfa_Control_Array(36));
    nfa_dfa_Control_Array37 <= std_logic_vector(tmp_nfa_dfa_Control_Array(37));
    nfa_dfa_Control_Array38 <= std_logic_vector(tmp_nfa_dfa_Control_Array(38));
    nfa_dfa_Control_Array39 <= std_logic_vector(tmp_nfa_dfa_Control_Array(39));
    nfa_dfa_Control_Array40 <= std_logic_vector(tmp_nfa_dfa_Control_Array(40));
    nfa_dfa_Control_Array41 <= std_logic_vector(tmp_nfa_dfa_Control_Array(41));
    nfa_dfa_Control_Array42 <= std_logic_vector(tmp_nfa_dfa_Control_Array(42));
    nfa_dfa_Control_Array43 <= std_logic_vector(tmp_nfa_dfa_Control_Array(43));
    nfa_dfa_Control_Array44 <= std_logic_vector(tmp_nfa_dfa_Control_Array(44));
    nfa_dfa_Control_Array45 <= std_logic_vector(tmp_nfa_dfa_Control_Array(45));
    nfa_dfa_Control_Array46 <= std_logic_vector(tmp_nfa_dfa_Control_Array(46));
    nfa_dfa_Control_Array47 <= std_logic_vector(tmp_nfa_dfa_Control_Array(47));
    nfa_dfa_Control_Array48 <= std_logic_vector(tmp_nfa_dfa_Control_Array(48));
    nfa_dfa_Control_Array49 <= std_logic_vector(tmp_nfa_dfa_Control_Array(49));
    nfa_dfa_Control_Array50 <= std_logic_vector(tmp_nfa_dfa_Control_Array(50));
    nfa_dfa_Control_Array51 <= std_logic_vector(tmp_nfa_dfa_Control_Array(51));
    nfa_dfa_Control_Array52 <= std_logic_vector(tmp_nfa_dfa_Control_Array(52));
    nfa_dfa_Control_Array53 <= std_logic_vector(tmp_nfa_dfa_Control_Array(53));
    nfa_dfa_Control_Array54 <= std_logic_vector(tmp_nfa_dfa_Control_Array(54));
    nfa_dfa_Control_Array55 <= std_logic_vector(tmp_nfa_dfa_Control_Array(55));
    nfa_dfa_Control_Array56 <= std_logic_vector(tmp_nfa_dfa_Control_Array(56));
    nfa_dfa_Control_Array57 <= std_logic_vector(tmp_nfa_dfa_Control_Array(57));
    nfa_dfa_Control_Array58 <= std_logic_vector(tmp_nfa_dfa_Control_Array(58));
    nfa_dfa_Control_Array59 <= std_logic_vector(tmp_nfa_dfa_Control_Array(59));
    nfa_dfa_Control_Array60 <= std_logic_vector(tmp_nfa_dfa_Control_Array(60));
    nfa_dfa_Control_Array61 <= std_logic_vector(tmp_nfa_dfa_Control_Array(61));
    nfa_dfa_Control_Array62 <= std_logic_vector(tmp_nfa_dfa_Control_Array(62));
    nfa_dfa_Control_Array63 <= std_logic_vector(tmp_nfa_dfa_Control_Array(63));
    nfa_dfa_Control_Array64 <= std_logic_vector(tmp_nfa_dfa_Control_Array(64));
    nfa_dfa_Control_Array65 <= std_logic_vector(tmp_nfa_dfa_Control_Array(65));
    nfa_dfa_Control_Array66 <= std_logic_vector(tmp_nfa_dfa_Control_Array(66));
    nfa_dfa_Control_Array67 <= std_logic_vector(tmp_nfa_dfa_Control_Array(67));
    nfa_dfa_Control_Array68 <= std_logic_vector(tmp_nfa_dfa_Control_Array(68));
    nfa_dfa_Control_Array69 <= std_logic_vector(tmp_nfa_dfa_Control_Array(69));
    nfa_dfa_Control_Array70 <= std_logic_vector(tmp_nfa_dfa_Control_Array(70));
    nfa_dfa_Control_Array71 <= std_logic_vector(tmp_nfa_dfa_Control_Array(71));
    nfa_dfa_Control_Array72 <= std_logic_vector(tmp_nfa_dfa_Control_Array(72));
    nfa_dfa_Control_Array73 <= std_logic_vector(tmp_nfa_dfa_Control_Array(73));
    nfa_dfa_Control_Array74 <= std_logic_vector(tmp_nfa_dfa_Control_Array(74));
    nfa_dfa_Control_Array75 <= std_logic_vector(tmp_nfa_dfa_Control_Array(75));
    nfa_dfa_Control_Array76 <= std_logic_vector(tmp_nfa_dfa_Control_Array(76));
    nfa_dfa_Control_Array77 <= std_logic_vector(tmp_nfa_dfa_Control_Array(77));
    nfa_dfa_Control_Array78 <= std_logic_vector(tmp_nfa_dfa_Control_Array(78));
    nfa_dfa_Control_Array79 <= std_logic_vector(tmp_nfa_dfa_Control_Array(79));
    nfa_dfa_Control_Array80 <= std_logic_vector(tmp_nfa_dfa_Control_Array(80));
    nfa_dfa_Control_Array81 <= std_logic_vector(tmp_nfa_dfa_Control_Array(81));
    nfa_dfa_Control_Array82 <= std_logic_vector(tmp_nfa_dfa_Control_Array(82));
    nfa_dfa_Control_Array83 <= std_logic_vector(tmp_nfa_dfa_Control_Array(83));
    nfa_dfa_Control_Array84 <= std_logic_vector(tmp_nfa_dfa_Control_Array(84));
    nfa_dfa_Control_Array85 <= std_logic_vector(tmp_nfa_dfa_Control_Array(85));
    nfa_dfa_Control_Array86 <= std_logic_vector(tmp_nfa_dfa_Control_Array(86));
    nfa_dfa_Control_Array87 <= std_logic_vector(tmp_nfa_dfa_Control_Array(87));
    nfa_dfa_Control_Array88 <= std_logic_vector(tmp_nfa_dfa_Control_Array(88));
    nfa_dfa_Control_Array89 <= std_logic_vector(tmp_nfa_dfa_Control_Array(89));
    nfa_dfa_Control_Array90 <= std_logic_vector(tmp_nfa_dfa_Control_Array(90));
    nfa_dfa_Control_Array91 <= std_logic_vector(tmp_nfa_dfa_Control_Array(91));
    nfa_dfa_Control_Array92 <= std_logic_vector(tmp_nfa_dfa_Control_Array(92));
    nfa_dfa_Control_Array93 <= std_logic_vector(tmp_nfa_dfa_Control_Array(93));
    nfa_dfa_Control_Array94 <= std_logic_vector(tmp_nfa_dfa_Control_Array(94));
    nfa_dfa_Control_Array95 <= std_logic_vector(tmp_nfa_dfa_Control_Array(95));
    nfa_dfa_Control_Array96 <= std_logic_vector(tmp_nfa_dfa_Control_Array(96));
    nfa_dfa_Control_Array97 <= std_logic_vector(tmp_nfa_dfa_Control_Array(97));
    nfa_dfa_Control_Array98 <= std_logic_vector(tmp_nfa_dfa_Control_Array(98));
    nfa_dfa_Control_Array99 <= std_logic_vector(tmp_nfa_dfa_Control_Array(99));
    nfa_dfa_Control_Array100 <= std_logic_vector(tmp_nfa_dfa_Control_Array(100));
    nfa_dfa_Control_Array101 <= std_logic_vector(tmp_nfa_dfa_Control_Array(101));
    nfa_dfa_Control_Array102 <= std_logic_vector(tmp_nfa_dfa_Control_Array(102));
    nfa_dfa_Control_Array103 <= std_logic_vector(tmp_nfa_dfa_Control_Array(103));
    nfa_dfa_Control_Array104 <= std_logic_vector(tmp_nfa_dfa_Control_Array(104));
    nfa_dfa_Control_Array105 <= std_logic_vector(tmp_nfa_dfa_Control_Array(105));
    nfa_dfa_Control_Array106 <= std_logic_vector(tmp_nfa_dfa_Control_Array(106));
    nfa_dfa_Control_Array107 <= std_logic_vector(tmp_nfa_dfa_Control_Array(107));
    nfa_dfa_Control_Array108 <= std_logic_vector(tmp_nfa_dfa_Control_Array(108));
    nfa_dfa_Control_Array109 <= std_logic_vector(tmp_nfa_dfa_Control_Array(109));
    nfa_dfa_Control_Array110 <= std_logic_vector(tmp_nfa_dfa_Control_Array(110));
    nfa_dfa_Control_Array111 <= std_logic_vector(tmp_nfa_dfa_Control_Array(111));
    nfa_dfa_Control_Array112 <= std_logic_vector(tmp_nfa_dfa_Control_Array(112));
    nfa_dfa_Control_Array113 <= std_logic_vector(tmp_nfa_dfa_Control_Array(113));
    nfa_dfa_Control_Array114 <= std_logic_vector(tmp_nfa_dfa_Control_Array(114));
    nfa_dfa_Control_Array115 <= std_logic_vector(tmp_nfa_dfa_Control_Array(115));
    nfa_dfa_Control_Array116 <= std_logic_vector(tmp_nfa_dfa_Control_Array(116));
    nfa_dfa_Control_Array117 <= std_logic_vector(tmp_nfa_dfa_Control_Array(117));
    nfa_dfa_Control_Array118 <= std_logic_vector(tmp_nfa_dfa_Control_Array(118));
    nfa_dfa_Control_Array119 <= std_logic_vector(tmp_nfa_dfa_Control_Array(119));
    nfa_dfa_Control_Array120 <= std_logic_vector(tmp_nfa_dfa_Control_Array(120));
    nfa_dfa_Control_Array121 <= std_logic_vector(tmp_nfa_dfa_Control_Array(121));
    nfa_dfa_Control_Array122 <= std_logic_vector(tmp_nfa_dfa_Control_Array(122));
    nfa_dfa_Control_Array123 <= std_logic_vector(tmp_nfa_dfa_Control_Array(123));
    nfa_dfa_Control_Array124 <= std_logic_vector(tmp_nfa_dfa_Control_Array(124));
    nfa_dfa_Control_Array125 <= std_logic_vector(tmp_nfa_dfa_Control_Array(125));
    nfa_dfa_Control_Array126 <= std_logic_vector(tmp_nfa_dfa_Control_Array(126));
    nfa_dfa_Control_Array127 <= std_logic_vector(tmp_nfa_dfa_Control_Array(127));
    nfa_dfa_Control_Array128 <= std_logic_vector(tmp_nfa_dfa_Control_Array(128));
    nfa_dfa_Control_Array129 <= std_logic_vector(tmp_nfa_dfa_Control_Array(129));
    nfa_dfa_Control_Array130 <= std_logic_vector(tmp_nfa_dfa_Control_Array(130));
    nfa_dfa_Control_Array131 <= std_logic_vector(tmp_nfa_dfa_Control_Array(131));
    nfa_dfa_Control_Array132 <= std_logic_vector(tmp_nfa_dfa_Control_Array(132));
    nfa_dfa_Control_Array133 <= std_logic_vector(tmp_nfa_dfa_Control_Array(133));
    nfa_dfa_Control_Array134 <= std_logic_vector(tmp_nfa_dfa_Control_Array(134));
    nfa_dfa_Control_Array135 <= std_logic_vector(tmp_nfa_dfa_Control_Array(135));
    nfa_dfa_Control_Array136 <= std_logic_vector(tmp_nfa_dfa_Control_Array(136));
    nfa_dfa_Control_Array137 <= std_logic_vector(tmp_nfa_dfa_Control_Array(137));
    nfa_dfa_Control_Array138 <= std_logic_vector(tmp_nfa_dfa_Control_Array(138));
    nfa_dfa_Control_Array139 <= std_logic_vector(tmp_nfa_dfa_Control_Array(139));
    nfa_dfa_Control_Array140 <= std_logic_vector(tmp_nfa_dfa_Control_Array(140));
    nfa_dfa_Control_Array141 <= std_logic_vector(tmp_nfa_dfa_Control_Array(141));
    nfa_dfa_Control_Array142 <= std_logic_vector(tmp_nfa_dfa_Control_Array(142));
    nfa_dfa_Control_Array143 <= std_logic_vector(tmp_nfa_dfa_Control_Array(143));
    nfa_dfa_Control_Array144 <= std_logic_vector(tmp_nfa_dfa_Control_Array(144));
    nfa_dfa_Control_Array145 <= std_logic_vector(tmp_nfa_dfa_Control_Array(145));
    nfa_dfa_Control_Array146 <= std_logic_vector(tmp_nfa_dfa_Control_Array(146));
    nfa_dfa_Control_Array147 <= std_logic_vector(tmp_nfa_dfa_Control_Array(147));
    nfa_dfa_Control_Array148 <= std_logic_vector(tmp_nfa_dfa_Control_Array(148));
    nfa_dfa_Control_Array149 <= std_logic_vector(tmp_nfa_dfa_Control_Array(149));
    nfa_dfa_Control_Array150 <= std_logic_vector(tmp_nfa_dfa_Control_Array(150));
    nfa_dfa_Control_Array151 <= std_logic_vector(tmp_nfa_dfa_Control_Array(151));
    nfa_dfa_Control_Array152 <= std_logic_vector(tmp_nfa_dfa_Control_Array(152));
    nfa_dfa_Control_Array153 <= std_logic_vector(tmp_nfa_dfa_Control_Array(153));
    nfa_dfa_Control_Array154 <= std_logic_vector(tmp_nfa_dfa_Control_Array(154));
    nfa_dfa_Control_Array155 <= std_logic_vector(tmp_nfa_dfa_Control_Array(155));
    nfa_dfa_Control_Array156 <= std_logic_vector(tmp_nfa_dfa_Control_Array(156));
    nfa_dfa_Control_Array157 <= std_logic_vector(tmp_nfa_dfa_Control_Array(157));
    nfa_dfa_Control_Array158 <= std_logic_vector(tmp_nfa_dfa_Control_Array(158));
    nfa_dfa_Control_Array159 <= std_logic_vector(tmp_nfa_dfa_Control_Array(159));
    nfa_dfa_Control_Array160 <= std_logic_vector(tmp_nfa_dfa_Control_Array(160));
    nfa_dfa_Control_Array161 <= std_logic_vector(tmp_nfa_dfa_Control_Array(161));
    nfa_dfa_Control_Array162 <= std_logic_vector(tmp_nfa_dfa_Control_Array(162));
    nfa_dfa_Control_Array163 <= std_logic_vector(tmp_nfa_dfa_Control_Array(163));
    nfa_dfa_Control_Array164 <= std_logic_vector(tmp_nfa_dfa_Control_Array(164));
    nfa_dfa_Control_Array165 <= std_logic_vector(tmp_nfa_dfa_Control_Array(165));
    nfa_dfa_Control_Array166 <= std_logic_vector(tmp_nfa_dfa_Control_Array(166));
    nfa_dfa_Control_Array167 <= std_logic_vector(tmp_nfa_dfa_Control_Array(167));
    nfa_dfa_Control_Array168 <= std_logic_vector(tmp_nfa_dfa_Control_Array(168));
    nfa_dfa_Control_Array169 <= std_logic_vector(tmp_nfa_dfa_Control_Array(169));
    nfa_dfa_Control_Array170 <= std_logic_vector(tmp_nfa_dfa_Control_Array(170));
    nfa_dfa_Control_Array171 <= std_logic_vector(tmp_nfa_dfa_Control_Array(171));
    nfa_dfa_Control_Array172 <= std_logic_vector(tmp_nfa_dfa_Control_Array(172));
    nfa_dfa_Control_Array173 <= std_logic_vector(tmp_nfa_dfa_Control_Array(173));
    nfa_dfa_Control_Array174 <= std_logic_vector(tmp_nfa_dfa_Control_Array(174));
    nfa_dfa_Control_Array175 <= std_logic_vector(tmp_nfa_dfa_Control_Array(175));
    nfa_dfa_Control_Array176 <= std_logic_vector(tmp_nfa_dfa_Control_Array(176));
    nfa_dfa_Control_Array177 <= std_logic_vector(tmp_nfa_dfa_Control_Array(177));
    nfa_dfa_Control_Array178 <= std_logic_vector(tmp_nfa_dfa_Control_Array(178));
    nfa_dfa_Control_Array179 <= std_logic_vector(tmp_nfa_dfa_Control_Array(179));
    nfa_dfa_Control_Array180 <= std_logic_vector(tmp_nfa_dfa_Control_Array(180));
    nfa_dfa_Control_Array181 <= std_logic_vector(tmp_nfa_dfa_Control_Array(181));
    nfa_dfa_Control_Array182 <= std_logic_vector(tmp_nfa_dfa_Control_Array(182));
    nfa_dfa_Control_Array183 <= std_logic_vector(tmp_nfa_dfa_Control_Array(183));
    nfa_dfa_Control_Array184 <= std_logic_vector(tmp_nfa_dfa_Control_Array(184));
    nfa_dfa_Control_Array185 <= std_logic_vector(tmp_nfa_dfa_Control_Array(185));
    nfa_dfa_Control_Array186 <= std_logic_vector(tmp_nfa_dfa_Control_Array(186));
    nfa_dfa_Control_Array187 <= std_logic_vector(tmp_nfa_dfa_Control_Array(187));
    nfa_dfa_Control_Array188 <= std_logic_vector(tmp_nfa_dfa_Control_Array(188));
    nfa_dfa_Control_Array189 <= std_logic_vector(tmp_nfa_dfa_Control_Array(189));
    nfa_dfa_Control_Array190 <= std_logic_vector(tmp_nfa_dfa_Control_Array(190));
    nfa_dfa_Control_Array191 <= std_logic_vector(tmp_nfa_dfa_Control_Array(191));
    nfa_dfa_Control_Array192 <= std_logic_vector(tmp_nfa_dfa_Control_Array(192));
    nfa_dfa_Control_Array193 <= std_logic_vector(tmp_nfa_dfa_Control_Array(193));
    nfa_dfa_Control_Array194 <= std_logic_vector(tmp_nfa_dfa_Control_Array(194));
    nfa_dfa_Control_Array195 <= std_logic_vector(tmp_nfa_dfa_Control_Array(195));
    nfa_dfa_Control_Array196 <= std_logic_vector(tmp_nfa_dfa_Control_Array(196));
    nfa_dfa_Control_Array197 <= std_logic_vector(tmp_nfa_dfa_Control_Array(197));
    nfa_dfa_Control_Array198 <= std_logic_vector(tmp_nfa_dfa_Control_Array(198));
    nfa_dfa_Control_Array199 <= std_logic_vector(tmp_nfa_dfa_Control_Array(199));
    nfa_dfa_Control_Array200 <= std_logic_vector(tmp_nfa_dfa_Control_Array(200));
    nfa_dfa_Control_Array201 <= std_logic_vector(tmp_nfa_dfa_Control_Array(201));
    nfa_dfa_Control_Array202 <= std_logic_vector(tmp_nfa_dfa_Control_Array(202));
    nfa_dfa_Control_Array203 <= std_logic_vector(tmp_nfa_dfa_Control_Array(203));
    nfa_dfa_Control_Array204 <= std_logic_vector(tmp_nfa_dfa_Control_Array(204));
    nfa_dfa_Control_Array205 <= std_logic_vector(tmp_nfa_dfa_Control_Array(205));
    nfa_dfa_Control_Array206 <= std_logic_vector(tmp_nfa_dfa_Control_Array(206));
    nfa_dfa_Control_Array207 <= std_logic_vector(tmp_nfa_dfa_Control_Array(207));
    nfa_dfa_Control_Array208 <= std_logic_vector(tmp_nfa_dfa_Control_Array(208));
    nfa_dfa_Control_Array209 <= std_logic_vector(tmp_nfa_dfa_Control_Array(209));
    nfa_dfa_Control_Array210 <= std_logic_vector(tmp_nfa_dfa_Control_Array(210));
    nfa_dfa_Control_Array211 <= std_logic_vector(tmp_nfa_dfa_Control_Array(211));
    nfa_dfa_Control_Array212 <= std_logic_vector(tmp_nfa_dfa_Control_Array(212));
    nfa_dfa_Control_Array213 <= std_logic_vector(tmp_nfa_dfa_Control_Array(213));
    nfa_dfa_Control_Array214 <= std_logic_vector(tmp_nfa_dfa_Control_Array(214));
    nfa_dfa_Control_Array215 <= std_logic_vector(tmp_nfa_dfa_Control_Array(215));
    nfa_dfa_Control_Array216 <= std_logic_vector(tmp_nfa_dfa_Control_Array(216));
    nfa_dfa_Control_Array217 <= std_logic_vector(tmp_nfa_dfa_Control_Array(217));
    nfa_dfa_Control_Array218 <= std_logic_vector(tmp_nfa_dfa_Control_Array(218));
    nfa_dfa_Control_Array219 <= std_logic_vector(tmp_nfa_dfa_Control_Array(219));
    nfa_dfa_Control_Array220 <= std_logic_vector(tmp_nfa_dfa_Control_Array(220));
    nfa_dfa_Control_Array221 <= std_logic_vector(tmp_nfa_dfa_Control_Array(221));
    nfa_dfa_Control_Array222 <= std_logic_vector(tmp_nfa_dfa_Control_Array(222));
    nfa_dfa_Control_Array223 <= std_logic_vector(tmp_nfa_dfa_Control_Array(223));
    nfa_dfa_Control_Array224 <= std_logic_vector(tmp_nfa_dfa_Control_Array(224));
    nfa_dfa_Control_Array225 <= std_logic_vector(tmp_nfa_dfa_Control_Array(225));
    nfa_dfa_Control_Array226 <= std_logic_vector(tmp_nfa_dfa_Control_Array(226));
    nfa_dfa_Control_Array227 <= std_logic_vector(tmp_nfa_dfa_Control_Array(227));
    nfa_dfa_Control_Array228 <= std_logic_vector(tmp_nfa_dfa_Control_Array(228));
    nfa_dfa_Control_Array229 <= std_logic_vector(tmp_nfa_dfa_Control_Array(229));
    nfa_dfa_Control_Array230 <= std_logic_vector(tmp_nfa_dfa_Control_Array(230));
    nfa_dfa_Control_Array231 <= std_logic_vector(tmp_nfa_dfa_Control_Array(231));
    nfa_dfa_Control_Array232 <= std_logic_vector(tmp_nfa_dfa_Control_Array(232));
    nfa_dfa_Control_Array233 <= std_logic_vector(tmp_nfa_dfa_Control_Array(233));
    nfa_dfa_Control_Array234 <= std_logic_vector(tmp_nfa_dfa_Control_Array(234));
    nfa_dfa_Control_Array235 <= std_logic_vector(tmp_nfa_dfa_Control_Array(235));
    nfa_dfa_Control_Array236 <= std_logic_vector(tmp_nfa_dfa_Control_Array(236));
    nfa_dfa_Control_Array237 <= std_logic_vector(tmp_nfa_dfa_Control_Array(237));
    nfa_dfa_Control_Array238 <= std_logic_vector(tmp_nfa_dfa_Control_Array(238));
    nfa_dfa_Control_Array239 <= std_logic_vector(tmp_nfa_dfa_Control_Array(239));
    nfa_dfa_Control_Array240 <= std_logic_vector(tmp_nfa_dfa_Control_Array(240));
    nfa_dfa_Control_Array241 <= std_logic_vector(tmp_nfa_dfa_Control_Array(241));
    nfa_dfa_Control_Array242 <= std_logic_vector(tmp_nfa_dfa_Control_Array(242));
    nfa_dfa_Control_Array243 <= std_logic_vector(tmp_nfa_dfa_Control_Array(243));
    nfa_dfa_Control_Array244 <= std_logic_vector(tmp_nfa_dfa_Control_Array(244));
    nfa_dfa_Control_Array245 <= std_logic_vector(tmp_nfa_dfa_Control_Array(245));
    nfa_dfa_Control_Array246 <= std_logic_vector(tmp_nfa_dfa_Control_Array(246));
    nfa_dfa_Control_Array247 <= std_logic_vector(tmp_nfa_dfa_Control_Array(247));
    nfa_dfa_Control_Array248 <= std_logic_vector(tmp_nfa_dfa_Control_Array(248));
    nfa_dfa_Control_Array249 <= std_logic_vector(tmp_nfa_dfa_Control_Array(249));
    nfa_dfa_Control_Array250 <= std_logic_vector(tmp_nfa_dfa_Control_Array(250));
    nfa_dfa_Control_Array251 <= std_logic_vector(tmp_nfa_dfa_Control_Array(251));
    nfa_dfa_Control_Array252 <= std_logic_vector(tmp_nfa_dfa_Control_Array(252));
    nfa_dfa_Control_Array253 <= std_logic_vector(tmp_nfa_dfa_Control_Array(253));
    nfa_dfa_Control_Array254 <= std_logic_vector(tmp_nfa_dfa_Control_Array(254));
    nfa_dfa_Control_Array255 <= std_logic_vector(tmp_nfa_dfa_Control_Array(255));
    nfa_dfa_Control_Array256 <= std_logic_vector(tmp_nfa_dfa_Control_Array(256));
    nfa_dfa_Control_Array257 <= std_logic_vector(tmp_nfa_dfa_Control_Array(257));
    nfa_dfa_Control_Array258 <= std_logic_vector(tmp_nfa_dfa_Control_Array(258));
    nfa_dfa_Control_Array259 <= std_logic_vector(tmp_nfa_dfa_Control_Array(259));
    nfa_dfa_Control_Array260 <= std_logic_vector(tmp_nfa_dfa_Control_Array(260));
    nfa_dfa_Control_Array261 <= std_logic_vector(tmp_nfa_dfa_Control_Array(261));
    nfa_dfa_Control_Array262 <= std_logic_vector(tmp_nfa_dfa_Control_Array(262));
    nfa_dfa_Control_Array263 <= std_logic_vector(tmp_nfa_dfa_Control_Array(263));
    nfa_dfa_Control_Array264 <= std_logic_vector(tmp_nfa_dfa_Control_Array(264));
    nfa_dfa_Control_Array265 <= std_logic_vector(tmp_nfa_dfa_Control_Array(265));
    nfa_dfa_Control_Array266 <= std_logic_vector(tmp_nfa_dfa_Control_Array(266));
    nfa_dfa_Control_Array267 <= std_logic_vector(tmp_nfa_dfa_Control_Array(267));
    nfa_dfa_Control_Array268 <= std_logic_vector(tmp_nfa_dfa_Control_Array(268));
    nfa_dfa_Control_Array269 <= std_logic_vector(tmp_nfa_dfa_Control_Array(269));
    nfa_dfa_Control_Array270 <= std_logic_vector(tmp_nfa_dfa_Control_Array(270));
    nfa_dfa_Control_Array271 <= std_logic_vector(tmp_nfa_dfa_Control_Array(271));
    nfa_dfa_Control_Array272 <= std_logic_vector(tmp_nfa_dfa_Control_Array(272));
    nfa_dfa_Control_Array273 <= std_logic_vector(tmp_nfa_dfa_Control_Array(273));
    nfa_dfa_Control_Array274 <= std_logic_vector(tmp_nfa_dfa_Control_Array(274));
    nfa_dfa_Control_Array275 <= std_logic_vector(tmp_nfa_dfa_Control_Array(275));
    nfa_dfa_Control_Array276 <= std_logic_vector(tmp_nfa_dfa_Control_Array(276));
    nfa_dfa_Control_Array277 <= std_logic_vector(tmp_nfa_dfa_Control_Array(277));
    nfa_dfa_Control_Array278 <= std_logic_vector(tmp_nfa_dfa_Control_Array(278));
    nfa_dfa_Control_Array279 <= std_logic_vector(tmp_nfa_dfa_Control_Array(279));
    nfa_dfa_Control_Array280 <= std_logic_vector(tmp_nfa_dfa_Control_Array(280));
    nfa_dfa_Control_Array281 <= std_logic_vector(tmp_nfa_dfa_Control_Array(281));
    nfa_dfa_Control_Array282 <= std_logic_vector(tmp_nfa_dfa_Control_Array(282));
    nfa_dfa_Control_Array283 <= std_logic_vector(tmp_nfa_dfa_Control_Array(283));
    nfa_dfa_Control_Array284 <= std_logic_vector(tmp_nfa_dfa_Control_Array(284));
    nfa_dfa_Control_Array285 <= std_logic_vector(tmp_nfa_dfa_Control_Array(285));
    nfa_dfa_Control_Array286 <= std_logic_vector(tmp_nfa_dfa_Control_Array(286));
    nfa_dfa_Control_Array287 <= std_logic_vector(tmp_nfa_dfa_Control_Array(287));
    nfa_dfa_Control_Array288 <= std_logic_vector(tmp_nfa_dfa_Control_Array(288));
    nfa_dfa_Control_Array289 <= std_logic_vector(tmp_nfa_dfa_Control_Array(289));
    nfa_dfa_Control_Array290 <= std_logic_vector(tmp_nfa_dfa_Control_Array(290));
    nfa_dfa_Control_Array291 <= std_logic_vector(tmp_nfa_dfa_Control_Array(291));
    nfa_dfa_Control_Array292 <= std_logic_vector(tmp_nfa_dfa_Control_Array(292));
    nfa_dfa_Control_Array293 <= std_logic_vector(tmp_nfa_dfa_Control_Array(293));
    nfa_dfa_Control_Array294 <= std_logic_vector(tmp_nfa_dfa_Control_Array(294));
    nfa_dfa_Control_Array295 <= std_logic_vector(tmp_nfa_dfa_Control_Array(295));
    nfa_dfa_Control_Array296 <= std_logic_vector(tmp_nfa_dfa_Control_Array(296));
    nfa_dfa_Control_Array297 <= std_logic_vector(tmp_nfa_dfa_Control_Array(297));
    nfa_dfa_Control_Array298 <= std_logic_vector(tmp_nfa_dfa_Control_Array(298));
    nfa_dfa_Control_Array299 <= std_logic_vector(tmp_nfa_dfa_Control_Array(299));
    nfa_dfa_Control_Array300 <= std_logic_vector(tmp_nfa_dfa_Control_Array(300));
    nfa_dfa_Control_Array301 <= std_logic_vector(tmp_nfa_dfa_Control_Array(301));
    nfa_dfa_Control_Array302 <= std_logic_vector(tmp_nfa_dfa_Control_Array(302));
    nfa_dfa_Control_Array303 <= std_logic_vector(tmp_nfa_dfa_Control_Array(303));
    nfa_dfa_Control_Array304 <= std_logic_vector(tmp_nfa_dfa_Control_Array(304));
    nfa_dfa_Control_Array305 <= std_logic_vector(tmp_nfa_dfa_Control_Array(305));
    nfa_dfa_Control_Array306 <= std_logic_vector(tmp_nfa_dfa_Control_Array(306));
    nfa_dfa_Control_Array307 <= std_logic_vector(tmp_nfa_dfa_Control_Array(307));
    nfa_dfa_Control_Array308 <= std_logic_vector(tmp_nfa_dfa_Control_Array(308));
    nfa_dfa_Control_Array309 <= std_logic_vector(tmp_nfa_dfa_Control_Array(309));
    nfa_dfa_Control_Array310 <= std_logic_vector(tmp_nfa_dfa_Control_Array(310));
    nfa_dfa_Control_Array311 <= std_logic_vector(tmp_nfa_dfa_Control_Array(311));
    nfa_dfa_Control_Array312 <= std_logic_vector(tmp_nfa_dfa_Control_Array(312));
    nfa_dfa_Control_Array313 <= std_logic_vector(tmp_nfa_dfa_Control_Array(313));
    nfa_dfa_Control_Array314 <= std_logic_vector(tmp_nfa_dfa_Control_Array(314));
    nfa_dfa_Control_Array315 <= std_logic_vector(tmp_nfa_dfa_Control_Array(315));
    nfa_dfa_Control_Array316 <= std_logic_vector(tmp_nfa_dfa_Control_Array(316));
    nfa_dfa_Control_Array317 <= std_logic_vector(tmp_nfa_dfa_Control_Array(317));
    nfa_dfa_Control_Array318 <= std_logic_vector(tmp_nfa_dfa_Control_Array(318));
    nfa_dfa_Control_Array319 <= std_logic_vector(tmp_nfa_dfa_Control_Array(319));
    nfa_dfa_Control_Array320 <= std_logic_vector(tmp_nfa_dfa_Control_Array(320));
    nfa_dfa_Control_Array321 <= std_logic_vector(tmp_nfa_dfa_Control_Array(321));
    nfa_dfa_Control_Array322 <= std_logic_vector(tmp_nfa_dfa_Control_Array(322));
    nfa_dfa_Control_Array323 <= std_logic_vector(tmp_nfa_dfa_Control_Array(323));
    nfa_dfa_Control_Array324 <= std_logic_vector(tmp_nfa_dfa_Control_Array(324));
    nfa_dfa_Control_Array325 <= std_logic_vector(tmp_nfa_dfa_Control_Array(325));
    nfa_dfa_Control_Array326 <= std_logic_vector(tmp_nfa_dfa_Control_Array(326));
    nfa_dfa_Control_Array327 <= std_logic_vector(tmp_nfa_dfa_Control_Array(327));
    nfa_dfa_Control_Array328 <= std_logic_vector(tmp_nfa_dfa_Control_Array(328));
    nfa_dfa_Control_Array329 <= std_logic_vector(tmp_nfa_dfa_Control_Array(329));
    nfa_dfa_Control_Array330 <= std_logic_vector(tmp_nfa_dfa_Control_Array(330));
    nfa_dfa_Control_Array331 <= std_logic_vector(tmp_nfa_dfa_Control_Array(331));
    nfa_dfa_Control_Array332 <= std_logic_vector(tmp_nfa_dfa_Control_Array(332));
    nfa_dfa_Control_Array333 <= std_logic_vector(tmp_nfa_dfa_Control_Array(333));
    nfa_dfa_Control_Array334 <= std_logic_vector(tmp_nfa_dfa_Control_Array(334));
    nfa_dfa_Control_Array335 <= std_logic_vector(tmp_nfa_dfa_Control_Array(335));
    nfa_dfa_Control_Array336 <= std_logic_vector(tmp_nfa_dfa_Control_Array(336));
    nfa_dfa_Control_Array337 <= std_logic_vector(tmp_nfa_dfa_Control_Array(337));
    nfa_dfa_Control_Array338 <= std_logic_vector(tmp_nfa_dfa_Control_Array(338));
    nfa_dfa_Control_Array339 <= std_logic_vector(tmp_nfa_dfa_Control_Array(339));
    nfa_dfa_Control_Array340 <= std_logic_vector(tmp_nfa_dfa_Control_Array(340));
    nfa_dfa_Control_Array341 <= std_logic_vector(tmp_nfa_dfa_Control_Array(341));
    nfa_dfa_Control_Array342 <= std_logic_vector(tmp_nfa_dfa_Control_Array(342));
    nfa_dfa_Control_Array343 <= std_logic_vector(tmp_nfa_dfa_Control_Array(343));
    nfa_dfa_Control_Array344 <= std_logic_vector(tmp_nfa_dfa_Control_Array(344));
    nfa_dfa_Control_Array345 <= std_logic_vector(tmp_nfa_dfa_Control_Array(345));
    nfa_dfa_Control_Array346 <= std_logic_vector(tmp_nfa_dfa_Control_Array(346));
    nfa_dfa_Control_Array347 <= std_logic_vector(tmp_nfa_dfa_Control_Array(347));
    nfa_dfa_Control_Array348 <= std_logic_vector(tmp_nfa_dfa_Control_Array(348));
    nfa_dfa_Control_Array349 <= std_logic_vector(tmp_nfa_dfa_Control_Array(349));
    nfa_dfa_Control_Array350 <= std_logic_vector(tmp_nfa_dfa_Control_Array(350));
    nfa_dfa_Control_Array351 <= std_logic_vector(tmp_nfa_dfa_Control_Array(351));
    nfa_dfa_Control_Array352 <= std_logic_vector(tmp_nfa_dfa_Control_Array(352));
    nfa_dfa_Control_Array353 <= std_logic_vector(tmp_nfa_dfa_Control_Array(353));
    nfa_dfa_Control_Array354 <= std_logic_vector(tmp_nfa_dfa_Control_Array(354));
    nfa_dfa_Control_Array355 <= std_logic_vector(tmp_nfa_dfa_Control_Array(355));
    nfa_dfa_Control_Array356 <= std_logic_vector(tmp_nfa_dfa_Control_Array(356));
    nfa_dfa_Control_Array357 <= std_logic_vector(tmp_nfa_dfa_Control_Array(357));
    nfa_dfa_Control_Array358 <= std_logic_vector(tmp_nfa_dfa_Control_Array(358));
    nfa_dfa_Control_Array359 <= std_logic_vector(tmp_nfa_dfa_Control_Array(359));
    nfa_dfa_Control_Array360 <= std_logic_vector(tmp_nfa_dfa_Control_Array(360));
    nfa_dfa_Control_Array361 <= std_logic_vector(tmp_nfa_dfa_Control_Array(361));
    nfa_dfa_Control_Array362 <= std_logic_vector(tmp_nfa_dfa_Control_Array(362));
    nfa_dfa_Control_Array363 <= std_logic_vector(tmp_nfa_dfa_Control_Array(363));
    nfa_dfa_Control_Array364 <= std_logic_vector(tmp_nfa_dfa_Control_Array(364));
    nfa_dfa_Control_Array365 <= std_logic_vector(tmp_nfa_dfa_Control_Array(365));
    nfa_dfa_Control_Array366 <= std_logic_vector(tmp_nfa_dfa_Control_Array(366));
    nfa_dfa_Control_Array367 <= std_logic_vector(tmp_nfa_dfa_Control_Array(367));
    nfa_dfa_Control_Array368 <= std_logic_vector(tmp_nfa_dfa_Control_Array(368));
    nfa_dfa_Control_Array369 <= std_logic_vector(tmp_nfa_dfa_Control_Array(369));
    nfa_dfa_Control_Array370 <= std_logic_vector(tmp_nfa_dfa_Control_Array(370));
    nfa_dfa_Control_Array371 <= std_logic_vector(tmp_nfa_dfa_Control_Array(371));
    nfa_dfa_Control_Array372 <= std_logic_vector(tmp_nfa_dfa_Control_Array(372));
    nfa_dfa_Control_Array373 <= std_logic_vector(tmp_nfa_dfa_Control_Array(373));
    nfa_dfa_Control_Array374 <= std_logic_vector(tmp_nfa_dfa_Control_Array(374));
    nfa_dfa_Control_Array375 <= std_logic_vector(tmp_nfa_dfa_Control_Array(375));
    nfa_dfa_Control_Array376 <= std_logic_vector(tmp_nfa_dfa_Control_Array(376));
    nfa_dfa_Control_Array377 <= std_logic_vector(tmp_nfa_dfa_Control_Array(377));
    nfa_dfa_Control_Array378 <= std_logic_vector(tmp_nfa_dfa_Control_Array(378));
    nfa_dfa_Control_Array379 <= std_logic_vector(tmp_nfa_dfa_Control_Array(379));
    nfa_dfa_Control_Array380 <= std_logic_vector(tmp_nfa_dfa_Control_Array(380));
    nfa_dfa_Control_Array381 <= std_logic_vector(tmp_nfa_dfa_Control_Array(381));
    nfa_dfa_Control_Array382 <= std_logic_vector(tmp_nfa_dfa_Control_Array(382));
    nfa_dfa_Control_Array383 <= std_logic_vector(tmp_nfa_dfa_Control_Array(383));
    nfa_dfa_Control_Array384 <= std_logic_vector(tmp_nfa_dfa_Control_Array(384));
    nfa_dfa_Control_Array385 <= std_logic_vector(tmp_nfa_dfa_Control_Array(385));
    nfa_dfa_Control_Array386 <= std_logic_vector(tmp_nfa_dfa_Control_Array(386));
    nfa_dfa_Control_Array387 <= std_logic_vector(tmp_nfa_dfa_Control_Array(387));
    nfa_dfa_Control_Array388 <= std_logic_vector(tmp_nfa_dfa_Control_Array(388));
    nfa_dfa_Control_Array389 <= std_logic_vector(tmp_nfa_dfa_Control_Array(389));
    nfa_dfa_Control_Array390 <= std_logic_vector(tmp_nfa_dfa_Control_Array(390));
    nfa_dfa_Control_Array391 <= std_logic_vector(tmp_nfa_dfa_Control_Array(391));
    nfa_dfa_Control_Array392 <= std_logic_vector(tmp_nfa_dfa_Control_Array(392));
    nfa_dfa_Control_Array393 <= std_logic_vector(tmp_nfa_dfa_Control_Array(393));
    nfa_dfa_Control_Array394 <= std_logic_vector(tmp_nfa_dfa_Control_Array(394));
    nfa_dfa_Control_Array395 <= std_logic_vector(tmp_nfa_dfa_Control_Array(395));
    nfa_dfa_Control_Array396 <= std_logic_vector(tmp_nfa_dfa_Control_Array(396));
    nfa_dfa_Control_Array397 <= std_logic_vector(tmp_nfa_dfa_Control_Array(397));
    nfa_dfa_Control_Array398 <= std_logic_vector(tmp_nfa_dfa_Control_Array(398));
    nfa_dfa_Control_Array399 <= std_logic_vector(tmp_nfa_dfa_Control_Array(399));
    nfa_dfa_Control_Array400 <= std_logic_vector(tmp_nfa_dfa_Control_Array(400));
    nfa_dfa_Control_Array401 <= std_logic_vector(tmp_nfa_dfa_Control_Array(401));
    nfa_dfa_Control_Array402 <= std_logic_vector(tmp_nfa_dfa_Control_Array(402));
    nfa_dfa_Control_Array403 <= std_logic_vector(tmp_nfa_dfa_Control_Array(403));
    nfa_dfa_Control_Array404 <= std_logic_vector(tmp_nfa_dfa_Control_Array(404));
    nfa_dfa_Control_Array405 <= std_logic_vector(tmp_nfa_dfa_Control_Array(405));
    nfa_dfa_Control_Array406 <= std_logic_vector(tmp_nfa_dfa_Control_Array(406));
    nfa_dfa_Control_Array407 <= std_logic_vector(tmp_nfa_dfa_Control_Array(407));
    nfa_dfa_Control_Array408 <= std_logic_vector(tmp_nfa_dfa_Control_Array(408));
    nfa_dfa_Control_Array409 <= std_logic_vector(tmp_nfa_dfa_Control_Array(409));
    nfa_dfa_Control_Array410 <= std_logic_vector(tmp_nfa_dfa_Control_Array(410));
    nfa_dfa_Control_Array411 <= std_logic_vector(tmp_nfa_dfa_Control_Array(411));
    nfa_dfa_Control_Array412 <= std_logic_vector(tmp_nfa_dfa_Control_Array(412));
    nfa_dfa_Control_Array413 <= std_logic_vector(tmp_nfa_dfa_Control_Array(413));
    nfa_dfa_Control_Array414 <= std_logic_vector(tmp_nfa_dfa_Control_Array(414));
    nfa_dfa_Control_Array415 <= std_logic_vector(tmp_nfa_dfa_Control_Array(415));
    nfa_dfa_Control_Array416 <= std_logic_vector(tmp_nfa_dfa_Control_Array(416));
    nfa_dfa_Control_Array417 <= std_logic_vector(tmp_nfa_dfa_Control_Array(417));
    nfa_dfa_Control_Array418 <= std_logic_vector(tmp_nfa_dfa_Control_Array(418));
    nfa_dfa_Control_Array419 <= std_logic_vector(tmp_nfa_dfa_Control_Array(419));
    nfa_dfa_Control_Array420 <= std_logic_vector(tmp_nfa_dfa_Control_Array(420));
    nfa_dfa_Control_Array421 <= std_logic_vector(tmp_nfa_dfa_Control_Array(421));
    nfa_dfa_Control_Array422 <= std_logic_vector(tmp_nfa_dfa_Control_Array(422));
    nfa_dfa_Control_Array423 <= std_logic_vector(tmp_nfa_dfa_Control_Array(423));
    nfa_dfa_Control_Array424 <= std_logic_vector(tmp_nfa_dfa_Control_Array(424));
    nfa_dfa_Control_Array425 <= std_logic_vector(tmp_nfa_dfa_Control_Array(425));
    nfa_dfa_Control_Array426 <= std_logic_vector(tmp_nfa_dfa_Control_Array(426));
    nfa_dfa_Control_Array427 <= std_logic_vector(tmp_nfa_dfa_Control_Array(427));
    nfa_dfa_Control_Array428 <= std_logic_vector(tmp_nfa_dfa_Control_Array(428));
    nfa_dfa_Control_Array429 <= std_logic_vector(tmp_nfa_dfa_Control_Array(429));
    nfa_dfa_Control_Array430 <= std_logic_vector(tmp_nfa_dfa_Control_Array(430));
    nfa_dfa_Control_Array431 <= std_logic_vector(tmp_nfa_dfa_Control_Array(431));
    nfa_dfa_Control_Array432 <= std_logic_vector(tmp_nfa_dfa_Control_Array(432));
    nfa_dfa_Control_Array433 <= std_logic_vector(tmp_nfa_dfa_Control_Array(433));
    nfa_dfa_Control_Array434 <= std_logic_vector(tmp_nfa_dfa_Control_Array(434));
    nfa_dfa_Control_Array435 <= std_logic_vector(tmp_nfa_dfa_Control_Array(435));
    nfa_dfa_Control_Array436 <= std_logic_vector(tmp_nfa_dfa_Control_Array(436));
    nfa_dfa_Control_Array437 <= std_logic_vector(tmp_nfa_dfa_Control_Array(437));
    nfa_dfa_Control_Array438 <= std_logic_vector(tmp_nfa_dfa_Control_Array(438));
    nfa_dfa_Control_Array439 <= std_logic_vector(tmp_nfa_dfa_Control_Array(439));
    nfa_dfa_Control_Array440 <= std_logic_vector(tmp_nfa_dfa_Control_Array(440));
    nfa_dfa_Control_Array441 <= std_logic_vector(tmp_nfa_dfa_Control_Array(441));
    nfa_dfa_Control_Array442 <= std_logic_vector(tmp_nfa_dfa_Control_Array(442));
    nfa_dfa_Control_Array443 <= std_logic_vector(tmp_nfa_dfa_Control_Array(443));
    nfa_dfa_Control_Array444 <= std_logic_vector(tmp_nfa_dfa_Control_Array(444));
    nfa_dfa_Control_Array445 <= std_logic_vector(tmp_nfa_dfa_Control_Array(445));
    nfa_dfa_Control_Array446 <= std_logic_vector(tmp_nfa_dfa_Control_Array(446));
    nfa_dfa_Control_Array447 <= std_logic_vector(tmp_nfa_dfa_Control_Array(447));
    nfa_dfa_Control_Array448 <= std_logic_vector(tmp_nfa_dfa_Control_Array(448));
    nfa_dfa_Control_Array449 <= std_logic_vector(tmp_nfa_dfa_Control_Array(449));
    nfa_dfa_Control_Array450 <= std_logic_vector(tmp_nfa_dfa_Control_Array(450));
    nfa_dfa_Control_Array451 <= std_logic_vector(tmp_nfa_dfa_Control_Array(451));
    nfa_dfa_Control_Array452 <= std_logic_vector(tmp_nfa_dfa_Control_Array(452));
    nfa_dfa_Control_Array453 <= std_logic_vector(tmp_nfa_dfa_Control_Array(453));
    nfa_dfa_Control_Array454 <= std_logic_vector(tmp_nfa_dfa_Control_Array(454));
    nfa_dfa_Control_Array455 <= std_logic_vector(tmp_nfa_dfa_Control_Array(455));
    nfa_dfa_Control_Array456 <= std_logic_vector(tmp_nfa_dfa_Control_Array(456));
    nfa_dfa_Control_Array457 <= std_logic_vector(tmp_nfa_dfa_Control_Array(457));
    nfa_dfa_Control_Array458 <= std_logic_vector(tmp_nfa_dfa_Control_Array(458));
    nfa_dfa_Control_Array459 <= std_logic_vector(tmp_nfa_dfa_Control_Array(459));
    nfa_dfa_Control_Array460 <= std_logic_vector(tmp_nfa_dfa_Control_Array(460));
    nfa_dfa_Control_Array461 <= std_logic_vector(tmp_nfa_dfa_Control_Array(461));
    nfa_dfa_Control_Array462 <= std_logic_vector(tmp_nfa_dfa_Control_Array(462));
    nfa_dfa_Control_Array463 <= std_logic_vector(tmp_nfa_dfa_Control_Array(463));
    nfa_dfa_Control_Array464 <= std_logic_vector(tmp_nfa_dfa_Control_Array(464));
    nfa_dfa_Control_Array465 <= std_logic_vector(tmp_nfa_dfa_Control_Array(465));
    nfa_dfa_Control_Array466 <= std_logic_vector(tmp_nfa_dfa_Control_Array(466));
    nfa_dfa_Control_Array467 <= std_logic_vector(tmp_nfa_dfa_Control_Array(467));
    nfa_dfa_Control_Array468 <= std_logic_vector(tmp_nfa_dfa_Control_Array(468));
    nfa_dfa_Control_Array469 <= std_logic_vector(tmp_nfa_dfa_Control_Array(469));
    nfa_dfa_Control_Array470 <= std_logic_vector(tmp_nfa_dfa_Control_Array(470));
    nfa_dfa_Control_Array471 <= std_logic_vector(tmp_nfa_dfa_Control_Array(471));
    nfa_dfa_Control_Array472 <= std_logic_vector(tmp_nfa_dfa_Control_Array(472));
    nfa_dfa_Control_Array473 <= std_logic_vector(tmp_nfa_dfa_Control_Array(473));
    nfa_dfa_Control_Array474 <= std_logic_vector(tmp_nfa_dfa_Control_Array(474));
    nfa_dfa_Control_Array475 <= std_logic_vector(tmp_nfa_dfa_Control_Array(475));
    nfa_dfa_Control_Array476 <= std_logic_vector(tmp_nfa_dfa_Control_Array(476));
    nfa_dfa_Control_Array477 <= std_logic_vector(tmp_nfa_dfa_Control_Array(477));
    nfa_dfa_Control_Array478 <= std_logic_vector(tmp_nfa_dfa_Control_Array(478));
    nfa_dfa_Control_Array479 <= std_logic_vector(tmp_nfa_dfa_Control_Array(479));
    nfa_dfa_Control_Array480 <= std_logic_vector(tmp_nfa_dfa_Control_Array(480));
    nfa_dfa_Control_Array481 <= std_logic_vector(tmp_nfa_dfa_Control_Array(481));
    nfa_dfa_Control_Array482 <= std_logic_vector(tmp_nfa_dfa_Control_Array(482));
    nfa_dfa_Control_Array483 <= std_logic_vector(tmp_nfa_dfa_Control_Array(483));
    nfa_dfa_Control_Array484 <= std_logic_vector(tmp_nfa_dfa_Control_Array(484));
    nfa_dfa_Control_Array485 <= std_logic_vector(tmp_nfa_dfa_Control_Array(485));
    nfa_dfa_Control_Array486 <= std_logic_vector(tmp_nfa_dfa_Control_Array(486));
    nfa_dfa_Control_Array487 <= std_logic_vector(tmp_nfa_dfa_Control_Array(487));
    nfa_dfa_Control_Array488 <= std_logic_vector(tmp_nfa_dfa_Control_Array(488));
    nfa_dfa_Control_Array489 <= std_logic_vector(tmp_nfa_dfa_Control_Array(489));
    nfa_dfa_Control_Array490 <= std_logic_vector(tmp_nfa_dfa_Control_Array(490));
    nfa_dfa_Control_Array491 <= std_logic_vector(tmp_nfa_dfa_Control_Array(491));
    nfa_dfa_Control_Array492 <= std_logic_vector(tmp_nfa_dfa_Control_Array(492));
    nfa_dfa_Control_Array493 <= std_logic_vector(tmp_nfa_dfa_Control_Array(493));
    nfa_dfa_Control_Array494 <= std_logic_vector(tmp_nfa_dfa_Control_Array(494));
    nfa_dfa_Control_Array495 <= std_logic_vector(tmp_nfa_dfa_Control_Array(495));
    nfa_dfa_Control_Array496 <= std_logic_vector(tmp_nfa_dfa_Control_Array(496));
    nfa_dfa_Control_Array497 <= std_logic_vector(tmp_nfa_dfa_Control_Array(497));
    nfa_dfa_Control_Array498 <= std_logic_vector(tmp_nfa_dfa_Control_Array(498));
    nfa_dfa_Control_Array499 <= std_logic_vector(tmp_nfa_dfa_Control_Array(499));
    nfa_dfa_Control_Array500 <= std_logic_vector(tmp_nfa_dfa_Control_Array(500));
    nfa_dfa_Control_Array501 <= std_logic_vector(tmp_nfa_dfa_Control_Array(501));
    nfa_dfa_Control_Array502 <= std_logic_vector(tmp_nfa_dfa_Control_Array(502));
    nfa_dfa_Control_Array503 <= std_logic_vector(tmp_nfa_dfa_Control_Array(503));
    nfa_dfa_Control_Array504 <= std_logic_vector(tmp_nfa_dfa_Control_Array(504));
    nfa_dfa_Control_Array505 <= std_logic_vector(tmp_nfa_dfa_Control_Array(505));
    nfa_dfa_Control_Array506 <= std_logic_vector(tmp_nfa_dfa_Control_Array(506));
    nfa_dfa_Control_Array507 <= std_logic_vector(tmp_nfa_dfa_Control_Array(507));
    nfa_dfa_Control_Array508 <= std_logic_vector(tmp_nfa_dfa_Control_Array(508));
    nfa_dfa_Control_Array509 <= std_logic_vector(tmp_nfa_dfa_Control_Array(509));
    nfa_dfa_Control_Array510 <= std_logic_vector(tmp_nfa_dfa_Control_Array(510));
    nfa_dfa_Control_Array511 <= std_logic_vector(tmp_nfa_dfa_Control_Array(511));
    nfa_dfa_Control_Array512 <= std_logic_vector(tmp_nfa_dfa_Control_Array(512));
    nfa_dfa_Control_Array513 <= std_logic_vector(tmp_nfa_dfa_Control_Array(513));
    nfa_dfa_Control_Array514 <= std_logic_vector(tmp_nfa_dfa_Control_Array(514));
    nfa_dfa_Control_Array515 <= std_logic_vector(tmp_nfa_dfa_Control_Array(515));
    nfa_dfa_Control_Array516 <= std_logic_vector(tmp_nfa_dfa_Control_Array(516));
    nfa_dfa_Control_Array517 <= std_logic_vector(tmp_nfa_dfa_Control_Array(517));
    nfa_dfa_Control_Array518 <= std_logic_vector(tmp_nfa_dfa_Control_Array(518));
    nfa_dfa_Control_Array519 <= std_logic_vector(tmp_nfa_dfa_Control_Array(519));
    nfa_dfa_Control_Array520 <= std_logic_vector(tmp_nfa_dfa_Control_Array(520));
    nfa_dfa_Control_Array521 <= std_logic_vector(tmp_nfa_dfa_Control_Array(521));
    nfa_dfa_Control_Array522 <= std_logic_vector(tmp_nfa_dfa_Control_Array(522));
    nfa_dfa_Control_Array523 <= std_logic_vector(tmp_nfa_dfa_Control_Array(523));
    nfa_dfa_Control_Array524 <= std_logic_vector(tmp_nfa_dfa_Control_Array(524));
    nfa_dfa_Control_Array525 <= std_logic_vector(tmp_nfa_dfa_Control_Array(525));
    nfa_dfa_Control_Array526 <= std_logic_vector(tmp_nfa_dfa_Control_Array(526));
    nfa_dfa_Control_Array527 <= std_logic_vector(tmp_nfa_dfa_Control_Array(527));
    nfa_dfa_Control_Array528 <= std_logic_vector(tmp_nfa_dfa_Control_Array(528));
    nfa_dfa_Control_Array529 <= std_logic_vector(tmp_nfa_dfa_Control_Array(529));
    nfa_dfa_Control_Array530 <= std_logic_vector(tmp_nfa_dfa_Control_Array(530));
    nfa_dfa_Control_Array531 <= std_logic_vector(tmp_nfa_dfa_Control_Array(531));
    nfa_dfa_Control_Array532 <= std_logic_vector(tmp_nfa_dfa_Control_Array(532));
    nfa_dfa_Control_Array533 <= std_logic_vector(tmp_nfa_dfa_Control_Array(533));
    nfa_dfa_Control_Array534 <= std_logic_vector(tmp_nfa_dfa_Control_Array(534));
    nfa_dfa_Control_Array535 <= std_logic_vector(tmp_nfa_dfa_Control_Array(535));
    nfa_dfa_Control_Array536 <= std_logic_vector(tmp_nfa_dfa_Control_Array(536));
    nfa_dfa_Control_Array537 <= std_logic_vector(tmp_nfa_dfa_Control_Array(537));
    nfa_dfa_Control_Array538 <= std_logic_vector(tmp_nfa_dfa_Control_Array(538));
    nfa_dfa_Control_Array539 <= std_logic_vector(tmp_nfa_dfa_Control_Array(539));
    nfa_dfa_Control_Array540 <= std_logic_vector(tmp_nfa_dfa_Control_Array(540));
    nfa_dfa_Control_Array541 <= std_logic_vector(tmp_nfa_dfa_Control_Array(541));
    nfa_dfa_Control_Array542 <= std_logic_vector(tmp_nfa_dfa_Control_Array(542));
    nfa_dfa_Control_Array543 <= std_logic_vector(tmp_nfa_dfa_Control_Array(543));
    nfa_dfa_Control_Array544 <= std_logic_vector(tmp_nfa_dfa_Control_Array(544));
    nfa_dfa_Control_Array545 <= std_logic_vector(tmp_nfa_dfa_Control_Array(545));
    nfa_dfa_Control_Array546 <= std_logic_vector(tmp_nfa_dfa_Control_Array(546));
    nfa_dfa_Control_Array547 <= std_logic_vector(tmp_nfa_dfa_Control_Array(547));
    nfa_dfa_Control_Array548 <= std_logic_vector(tmp_nfa_dfa_Control_Array(548));
    nfa_dfa_Control_Array549 <= std_logic_vector(tmp_nfa_dfa_Control_Array(549));
    nfa_dfa_Control_Array550 <= std_logic_vector(tmp_nfa_dfa_Control_Array(550));
    nfa_dfa_Control_Array551 <= std_logic_vector(tmp_nfa_dfa_Control_Array(551));
    nfa_dfa_Control_Array552 <= std_logic_vector(tmp_nfa_dfa_Control_Array(552));
    nfa_dfa_Control_Array553 <= std_logic_vector(tmp_nfa_dfa_Control_Array(553));
    nfa_dfa_Control_Array554 <= std_logic_vector(tmp_nfa_dfa_Control_Array(554));
    nfa_dfa_Control_Array555 <= std_logic_vector(tmp_nfa_dfa_Control_Array(555));
    nfa_dfa_Control_Array556 <= std_logic_vector(tmp_nfa_dfa_Control_Array(556));
    nfa_dfa_Control_Array557 <= std_logic_vector(tmp_nfa_dfa_Control_Array(557));
    nfa_dfa_Control_Array558 <= std_logic_vector(tmp_nfa_dfa_Control_Array(558));
    nfa_dfa_Control_Array559 <= std_logic_vector(tmp_nfa_dfa_Control_Array(559));
    nfa_dfa_Control_Array560 <= std_logic_vector(tmp_nfa_dfa_Control_Array(560));
    nfa_dfa_Control_Array561 <= std_logic_vector(tmp_nfa_dfa_Control_Array(561));
    nfa_dfa_Control_Array562 <= std_logic_vector(tmp_nfa_dfa_Control_Array(562));
    nfa_dfa_Control_Array563 <= std_logic_vector(tmp_nfa_dfa_Control_Array(563));
    nfa_dfa_Control_Array564 <= std_logic_vector(tmp_nfa_dfa_Control_Array(564));
    nfa_dfa_Control_Array565 <= std_logic_vector(tmp_nfa_dfa_Control_Array(565));
    nfa_dfa_Control_Array566 <= std_logic_vector(tmp_nfa_dfa_Control_Array(566));
    nfa_dfa_Control_Array567 <= std_logic_vector(tmp_nfa_dfa_Control_Array(567));
    nfa_dfa_Control_Array568 <= std_logic_vector(tmp_nfa_dfa_Control_Array(568));
    nfa_dfa_Control_Array569 <= std_logic_vector(tmp_nfa_dfa_Control_Array(569));
    nfa_dfa_Control_Array570 <= std_logic_vector(tmp_nfa_dfa_Control_Array(570));
    nfa_dfa_Control_Array571 <= std_logic_vector(tmp_nfa_dfa_Control_Array(571));
    nfa_dfa_Control_Array572 <= std_logic_vector(tmp_nfa_dfa_Control_Array(572));
    nfa_dfa_Control_Array573 <= std_logic_vector(tmp_nfa_dfa_Control_Array(573));
    nfa_dfa_Control_Array574 <= std_logic_vector(tmp_nfa_dfa_Control_Array(574));
    nfa_dfa_Control_Array575 <= std_logic_vector(tmp_nfa_dfa_Control_Array(575));
    nfa_dfa_Control_Array576 <= std_logic_vector(tmp_nfa_dfa_Control_Array(576));
    nfa_dfa_Control_Array577 <= std_logic_vector(tmp_nfa_dfa_Control_Array(577));
    nfa_dfa_Control_Array578 <= std_logic_vector(tmp_nfa_dfa_Control_Array(578));
    nfa_dfa_Control_Array579 <= std_logic_vector(tmp_nfa_dfa_Control_Array(579));
    nfa_dfa_Control_Array580 <= std_logic_vector(tmp_nfa_dfa_Control_Array(580));
    nfa_dfa_Control_Array581 <= std_logic_vector(tmp_nfa_dfa_Control_Array(581));
    nfa_dfa_Control_Array582 <= std_logic_vector(tmp_nfa_dfa_Control_Array(582));
    nfa_dfa_Control_Array583 <= std_logic_vector(tmp_nfa_dfa_Control_Array(583));
    nfa_dfa_Control_Array584 <= std_logic_vector(tmp_nfa_dfa_Control_Array(584));
    nfa_dfa_Control_Array585 <= std_logic_vector(tmp_nfa_dfa_Control_Array(585));
    nfa_dfa_Control_Array586 <= std_logic_vector(tmp_nfa_dfa_Control_Array(586));
    nfa_dfa_Control_Array587 <= std_logic_vector(tmp_nfa_dfa_Control_Array(587));
    nfa_dfa_Control_Array588 <= std_logic_vector(tmp_nfa_dfa_Control_Array(588));
    nfa_dfa_Control_Array589 <= std_logic_vector(tmp_nfa_dfa_Control_Array(589));
    nfa_dfa_Control_Array590 <= std_logic_vector(tmp_nfa_dfa_Control_Array(590));
    nfa_dfa_Control_Array591 <= std_logic_vector(tmp_nfa_dfa_Control_Array(591));
    nfa_dfa_Control_Array592 <= std_logic_vector(tmp_nfa_dfa_Control_Array(592));
    nfa_dfa_Control_Array593 <= std_logic_vector(tmp_nfa_dfa_Control_Array(593));
    nfa_dfa_Control_Array594 <= std_logic_vector(tmp_nfa_dfa_Control_Array(594));
    nfa_dfa_Control_Array595 <= std_logic_vector(tmp_nfa_dfa_Control_Array(595));
    nfa_dfa_Control_Array596 <= std_logic_vector(tmp_nfa_dfa_Control_Array(596));
    nfa_dfa_Control_Array597 <= std_logic_vector(tmp_nfa_dfa_Control_Array(597));
    nfa_dfa_Control_Array598 <= std_logic_vector(tmp_nfa_dfa_Control_Array(598));
    nfa_dfa_Control_Array599 <= std_logic_vector(tmp_nfa_dfa_Control_Array(599));
    nfa_dfa_Control_Array600 <= std_logic_vector(tmp_nfa_dfa_Control_Array(600));
    nfa_dfa_Control_Array601 <= std_logic_vector(tmp_nfa_dfa_Control_Array(601));
    nfa_dfa_Control_Array602 <= std_logic_vector(tmp_nfa_dfa_Control_Array(602));
    nfa_dfa_Control_Array603 <= std_logic_vector(tmp_nfa_dfa_Control_Array(603));
    nfa_dfa_Control_Array604 <= std_logic_vector(tmp_nfa_dfa_Control_Array(604));
    nfa_dfa_Control_Array605 <= std_logic_vector(tmp_nfa_dfa_Control_Array(605));
    nfa_dfa_Control_Array606 <= std_logic_vector(tmp_nfa_dfa_Control_Array(606));
    nfa_dfa_Control_Array607 <= std_logic_vector(tmp_nfa_dfa_Control_Array(607));
    nfa_dfa_Control_Array608 <= std_logic_vector(tmp_nfa_dfa_Control_Array(608));
    nfa_dfa_Control_Array609 <= std_logic_vector(tmp_nfa_dfa_Control_Array(609));
    nfa_dfa_Control_Array610 <= std_logic_vector(tmp_nfa_dfa_Control_Array(610));
    nfa_dfa_Control_Array611 <= std_logic_vector(tmp_nfa_dfa_Control_Array(611));
    nfa_dfa_Control_Array612 <= std_logic_vector(tmp_nfa_dfa_Control_Array(612));
    nfa_dfa_Control_Array613 <= std_logic_vector(tmp_nfa_dfa_Control_Array(613));
    nfa_dfa_Control_Array614 <= std_logic_vector(tmp_nfa_dfa_Control_Array(614));
    nfa_dfa_Control_Array615 <= std_logic_vector(tmp_nfa_dfa_Control_Array(615));
    nfa_dfa_Control_Array616 <= std_logic_vector(tmp_nfa_dfa_Control_Array(616));
    nfa_dfa_Control_Array617 <= std_logic_vector(tmp_nfa_dfa_Control_Array(617));
    nfa_dfa_Control_Array618 <= std_logic_vector(tmp_nfa_dfa_Control_Array(618));
    nfa_dfa_Control_Array619 <= std_logic_vector(tmp_nfa_dfa_Control_Array(619));
    nfa_dfa_Control_Array620 <= std_logic_vector(tmp_nfa_dfa_Control_Array(620));
    nfa_dfa_Control_Array621 <= std_logic_vector(tmp_nfa_dfa_Control_Array(621));
    nfa_dfa_Control_Array622 <= std_logic_vector(tmp_nfa_dfa_Control_Array(622));
    nfa_dfa_Control_Array623 <= std_logic_vector(tmp_nfa_dfa_Control_Array(623));
    nfa_dfa_Control_Array624 <= std_logic_vector(tmp_nfa_dfa_Control_Array(624));
    nfa_dfa_Control_Array625 <= std_logic_vector(tmp_nfa_dfa_Control_Array(625));
    nfa_dfa_Control_Array626 <= std_logic_vector(tmp_nfa_dfa_Control_Array(626));
    nfa_dfa_Control_Array627 <= std_logic_vector(tmp_nfa_dfa_Control_Array(627));
    nfa_dfa_Control_Array628 <= std_logic_vector(tmp_nfa_dfa_Control_Array(628));
    nfa_dfa_Control_Array629 <= std_logic_vector(tmp_nfa_dfa_Control_Array(629));
    nfa_dfa_Control_Array630 <= std_logic_vector(tmp_nfa_dfa_Control_Array(630));
    nfa_dfa_Control_Array631 <= std_logic_vector(tmp_nfa_dfa_Control_Array(631));
    nfa_dfa_Control_Array632 <= std_logic_vector(tmp_nfa_dfa_Control_Array(632));
    nfa_dfa_Control_Array633 <= std_logic_vector(tmp_nfa_dfa_Control_Array(633));
    nfa_dfa_Control_Array634 <= std_logic_vector(tmp_nfa_dfa_Control_Array(634));
    nfa_dfa_Control_Array635 <= std_logic_vector(tmp_nfa_dfa_Control_Array(635));
    nfa_dfa_Control_Array636 <= std_logic_vector(tmp_nfa_dfa_Control_Array(636));
    nfa_dfa_Control_Array637 <= std_logic_vector(tmp_nfa_dfa_Control_Array(637));
    nfa_dfa_Control_Array638 <= std_logic_vector(tmp_nfa_dfa_Control_Array(638));
    nfa_dfa_Control_Array639 <= std_logic_vector(tmp_nfa_dfa_Control_Array(639));
    nfa_dfa_Control_Array640 <= std_logic_vector(tmp_nfa_dfa_Control_Array(640));
    nfa_dfa_Control_Array641 <= std_logic_vector(tmp_nfa_dfa_Control_Array(641));
    nfa_dfa_Control_Array642 <= std_logic_vector(tmp_nfa_dfa_Control_Array(642));
    nfa_dfa_Control_Array643 <= std_logic_vector(tmp_nfa_dfa_Control_Array(643));
    nfa_dfa_Control_Array644 <= std_logic_vector(tmp_nfa_dfa_Control_Array(644));
    nfa_dfa_Control_Array645 <= std_logic_vector(tmp_nfa_dfa_Control_Array(645));
    nfa_dfa_Control_Array646 <= std_logic_vector(tmp_nfa_dfa_Control_Array(646));
    nfa_dfa_Control_Array647 <= std_logic_vector(tmp_nfa_dfa_Control_Array(647));
    nfa_dfa_Control_Array648 <= std_logic_vector(tmp_nfa_dfa_Control_Array(648));
    nfa_dfa_Control_Array649 <= std_logic_vector(tmp_nfa_dfa_Control_Array(649));
    nfa_dfa_Control_Array650 <= std_logic_vector(tmp_nfa_dfa_Control_Array(650));
    nfa_dfa_Control_Array651 <= std_logic_vector(tmp_nfa_dfa_Control_Array(651));
    nfa_dfa_Control_Array652 <= std_logic_vector(tmp_nfa_dfa_Control_Array(652));
    nfa_dfa_Control_Array653 <= std_logic_vector(tmp_nfa_dfa_Control_Array(653));
    nfa_dfa_Control_Array654 <= std_logic_vector(tmp_nfa_dfa_Control_Array(654));
    nfa_dfa_Control_Array655 <= std_logic_vector(tmp_nfa_dfa_Control_Array(655));
    nfa_dfa_Control_Array656 <= std_logic_vector(tmp_nfa_dfa_Control_Array(656));
    nfa_dfa_Control_Array657 <= std_logic_vector(tmp_nfa_dfa_Control_Array(657));
    nfa_dfa_Control_Array658 <= std_logic_vector(tmp_nfa_dfa_Control_Array(658));
    nfa_dfa_Control_Array659 <= std_logic_vector(tmp_nfa_dfa_Control_Array(659));
    nfa_dfa_Control_Array660 <= std_logic_vector(tmp_nfa_dfa_Control_Array(660));
    nfa_dfa_Control_Array661 <= std_logic_vector(tmp_nfa_dfa_Control_Array(661));
    nfa_dfa_Control_Array662 <= std_logic_vector(tmp_nfa_dfa_Control_Array(662));
    nfa_dfa_Control_Array663 <= std_logic_vector(tmp_nfa_dfa_Control_Array(663));
    nfa_dfa_Control_Array664 <= std_logic_vector(tmp_nfa_dfa_Control_Array(664));
    nfa_dfa_Control_Array665 <= std_logic_vector(tmp_nfa_dfa_Control_Array(665));
    nfa_dfa_Control_Array666 <= std_logic_vector(tmp_nfa_dfa_Control_Array(666));
    nfa_dfa_Control_Array667 <= std_logic_vector(tmp_nfa_dfa_Control_Array(667));
    nfa_dfa_Control_Array668 <= std_logic_vector(tmp_nfa_dfa_Control_Array(668));
    nfa_dfa_Control_Array669 <= std_logic_vector(tmp_nfa_dfa_Control_Array(669));
    nfa_dfa_Control_Array670 <= std_logic_vector(tmp_nfa_dfa_Control_Array(670));
    nfa_dfa_Control_Array671 <= std_logic_vector(tmp_nfa_dfa_Control_Array(671));
    nfa_dfa_Control_Array672 <= std_logic_vector(tmp_nfa_dfa_Control_Array(672));
    nfa_dfa_Control_Array673 <= std_logic_vector(tmp_nfa_dfa_Control_Array(673));
    nfa_dfa_Control_Array674 <= std_logic_vector(tmp_nfa_dfa_Control_Array(674));
    nfa_dfa_Control_Array675 <= std_logic_vector(tmp_nfa_dfa_Control_Array(675));
    nfa_dfa_Control_Array676 <= std_logic_vector(tmp_nfa_dfa_Control_Array(676));
    nfa_dfa_Control_Array677 <= std_logic_vector(tmp_nfa_dfa_Control_Array(677));
    nfa_dfa_Control_Array678 <= std_logic_vector(tmp_nfa_dfa_Control_Array(678));
    nfa_dfa_Control_Array679 <= std_logic_vector(tmp_nfa_dfa_Control_Array(679));
    nfa_dfa_Control_Array680 <= std_logic_vector(tmp_nfa_dfa_Control_Array(680));
    nfa_dfa_Control_Array681 <= std_logic_vector(tmp_nfa_dfa_Control_Array(681));
    nfa_dfa_Control_Array682 <= std_logic_vector(tmp_nfa_dfa_Control_Array(682));
    nfa_dfa_Control_Array683 <= std_logic_vector(tmp_nfa_dfa_Control_Array(683));
    nfa_dfa_Control_Array684 <= std_logic_vector(tmp_nfa_dfa_Control_Array(684));
    nfa_dfa_Control_Array685 <= std_logic_vector(tmp_nfa_dfa_Control_Array(685));
    nfa_dfa_Control_Array686 <= std_logic_vector(tmp_nfa_dfa_Control_Array(686));
    nfa_dfa_Control_Array687 <= std_logic_vector(tmp_nfa_dfa_Control_Array(687));
    nfa_dfa_Control_Array688 <= std_logic_vector(tmp_nfa_dfa_Control_Array(688));
    nfa_dfa_Control_Array689 <= std_logic_vector(tmp_nfa_dfa_Control_Array(689));
    nfa_dfa_Control_Array690 <= std_logic_vector(tmp_nfa_dfa_Control_Array(690));
    nfa_dfa_Control_Array691 <= std_logic_vector(tmp_nfa_dfa_Control_Array(691));
    nfa_dfa_Control_Array692 <= std_logic_vector(tmp_nfa_dfa_Control_Array(692));
    nfa_dfa_Control_Array693 <= std_logic_vector(tmp_nfa_dfa_Control_Array(693));
    nfa_dfa_Control_Array694 <= std_logic_vector(tmp_nfa_dfa_Control_Array(694));
    nfa_dfa_Control_Array695 <= std_logic_vector(tmp_nfa_dfa_Control_Array(695));
    nfa_dfa_Control_Array696 <= std_logic_vector(tmp_nfa_dfa_Control_Array(696));
    nfa_dfa_Control_Array697 <= std_logic_vector(tmp_nfa_dfa_Control_Array(697));
    nfa_dfa_Control_Array698 <= std_logic_vector(tmp_nfa_dfa_Control_Array(698));
    nfa_dfa_Control_Array699 <= std_logic_vector(tmp_nfa_dfa_Control_Array(699));
    nfa_dfa_Control_Array700 <= std_logic_vector(tmp_nfa_dfa_Control_Array(700));
    nfa_dfa_Control_Array701 <= std_logic_vector(tmp_nfa_dfa_Control_Array(701));
    nfa_dfa_Control_Array702 <= std_logic_vector(tmp_nfa_dfa_Control_Array(702));
    nfa_dfa_Control_Array703 <= std_logic_vector(tmp_nfa_dfa_Control_Array(703));
    nfa_dfa_Control_Array704 <= std_logic_vector(tmp_nfa_dfa_Control_Array(704));
    nfa_dfa_Control_Array705 <= std_logic_vector(tmp_nfa_dfa_Control_Array(705));
    nfa_dfa_Control_Array706 <= std_logic_vector(tmp_nfa_dfa_Control_Array(706));
    nfa_dfa_Control_Array707 <= std_logic_vector(tmp_nfa_dfa_Control_Array(707));
    nfa_dfa_Control_Array708 <= std_logic_vector(tmp_nfa_dfa_Control_Array(708));
    nfa_dfa_Control_Array709 <= std_logic_vector(tmp_nfa_dfa_Control_Array(709));
    nfa_dfa_Control_Array710 <= std_logic_vector(tmp_nfa_dfa_Control_Array(710));
    nfa_dfa_Control_Array711 <= std_logic_vector(tmp_nfa_dfa_Control_Array(711));
    nfa_dfa_Control_Array712 <= std_logic_vector(tmp_nfa_dfa_Control_Array(712));
    nfa_dfa_Control_Array713 <= std_logic_vector(tmp_nfa_dfa_Control_Array(713));
    nfa_dfa_Control_Array714 <= std_logic_vector(tmp_nfa_dfa_Control_Array(714));
    nfa_dfa_Control_Array715 <= std_logic_vector(tmp_nfa_dfa_Control_Array(715));
    nfa_dfa_Control_Array716 <= std_logic_vector(tmp_nfa_dfa_Control_Array(716));
    nfa_dfa_Control_Array717 <= std_logic_vector(tmp_nfa_dfa_Control_Array(717));
    nfa_dfa_Control_Array718 <= std_logic_vector(tmp_nfa_dfa_Control_Array(718));
    nfa_dfa_Control_Array719 <= std_logic_vector(tmp_nfa_dfa_Control_Array(719));
    nfa_dfa_Control_Array720 <= std_logic_vector(tmp_nfa_dfa_Control_Array(720));
    nfa_dfa_Control_Array721 <= std_logic_vector(tmp_nfa_dfa_Control_Array(721));
    nfa_dfa_Control_Array722 <= std_logic_vector(tmp_nfa_dfa_Control_Array(722));
    nfa_dfa_Control_Array723 <= std_logic_vector(tmp_nfa_dfa_Control_Array(723));
    nfa_dfa_Control_Array724 <= std_logic_vector(tmp_nfa_dfa_Control_Array(724));
    nfa_dfa_Control_Array725 <= std_logic_vector(tmp_nfa_dfa_Control_Array(725));
    nfa_dfa_Control_Array726 <= std_logic_vector(tmp_nfa_dfa_Control_Array(726));
    nfa_dfa_Control_Array727 <= std_logic_vector(tmp_nfa_dfa_Control_Array(727));
    nfa_dfa_Control_Array728 <= std_logic_vector(tmp_nfa_dfa_Control_Array(728));
    nfa_dfa_Control_Array729 <= std_logic_vector(tmp_nfa_dfa_Control_Array(729));
    nfa_dfa_Control_Array730 <= std_logic_vector(tmp_nfa_dfa_Control_Array(730));
    nfa_dfa_Control_Array731 <= std_logic_vector(tmp_nfa_dfa_Control_Array(731));
    nfa_dfa_Control_Array732 <= std_logic_vector(tmp_nfa_dfa_Control_Array(732));
    nfa_dfa_Control_Array733 <= std_logic_vector(tmp_nfa_dfa_Control_Array(733));
    nfa_dfa_Control_Array734 <= std_logic_vector(tmp_nfa_dfa_Control_Array(734));
    nfa_dfa_Control_Array735 <= std_logic_vector(tmp_nfa_dfa_Control_Array(735));
    nfa_dfa_Control_Array736 <= std_logic_vector(tmp_nfa_dfa_Control_Array(736));
    nfa_dfa_Control_Array737 <= std_logic_vector(tmp_nfa_dfa_Control_Array(737));
    nfa_dfa_Control_Array738 <= std_logic_vector(tmp_nfa_dfa_Control_Array(738));
    nfa_dfa_Control_Array739 <= std_logic_vector(tmp_nfa_dfa_Control_Array(739));
    nfa_dfa_Control_Array740 <= std_logic_vector(tmp_nfa_dfa_Control_Array(740));
    nfa_dfa_Control_Array741 <= std_logic_vector(tmp_nfa_dfa_Control_Array(741));
    nfa_dfa_Control_Array742 <= std_logic_vector(tmp_nfa_dfa_Control_Array(742));
    nfa_dfa_Control_Array743 <= std_logic_vector(tmp_nfa_dfa_Control_Array(743));
    nfa_dfa_Control_Array744 <= std_logic_vector(tmp_nfa_dfa_Control_Array(744));
    nfa_dfa_Control_Array745 <= std_logic_vector(tmp_nfa_dfa_Control_Array(745));
    nfa_dfa_Control_Array746 <= std_logic_vector(tmp_nfa_dfa_Control_Array(746));
    nfa_dfa_Control_Array747 <= std_logic_vector(tmp_nfa_dfa_Control_Array(747));
    nfa_dfa_Control_Array748 <= std_logic_vector(tmp_nfa_dfa_Control_Array(748));
    nfa_dfa_Control_Array749 <= std_logic_vector(tmp_nfa_dfa_Control_Array(749));
    nfa_dfa_Control_Array750 <= std_logic_vector(tmp_nfa_dfa_Control_Array(750));
    nfa_dfa_Control_Array751 <= std_logic_vector(tmp_nfa_dfa_Control_Array(751));
    nfa_dfa_Control_Array752 <= std_logic_vector(tmp_nfa_dfa_Control_Array(752));
    nfa_dfa_Control_Array753 <= std_logic_vector(tmp_nfa_dfa_Control_Array(753));
    nfa_dfa_Control_Array754 <= std_logic_vector(tmp_nfa_dfa_Control_Array(754));
    nfa_dfa_Control_Array755 <= std_logic_vector(tmp_nfa_dfa_Control_Array(755));
    nfa_dfa_Control_Array756 <= std_logic_vector(tmp_nfa_dfa_Control_Array(756));
    nfa_dfa_Control_Array757 <= std_logic_vector(tmp_nfa_dfa_Control_Array(757));
    nfa_dfa_Control_Array758 <= std_logic_vector(tmp_nfa_dfa_Control_Array(758));
    nfa_dfa_Control_Array759 <= std_logic_vector(tmp_nfa_dfa_Control_Array(759));
    nfa_dfa_Control_Array760 <= std_logic_vector(tmp_nfa_dfa_Control_Array(760));
    nfa_dfa_Control_Array761 <= std_logic_vector(tmp_nfa_dfa_Control_Array(761));
    nfa_dfa_Control_Array762 <= std_logic_vector(tmp_nfa_dfa_Control_Array(762));
    nfa_dfa_Control_Array763 <= std_logic_vector(tmp_nfa_dfa_Control_Array(763));
    nfa_dfa_Control_Array764 <= std_logic_vector(tmp_nfa_dfa_Control_Array(764));
    nfa_dfa_Control_Array765 <= std_logic_vector(tmp_nfa_dfa_Control_Array(765));
    nfa_dfa_Control_Array766 <= std_logic_vector(tmp_nfa_dfa_Control_Array(766));
    nfa_dfa_Control_Array767 <= std_logic_vector(tmp_nfa_dfa_Control_Array(767));
    nfa_dfa_Control_Array768 <= std_logic_vector(tmp_nfa_dfa_Control_Array(768));
    nfa_dfa_Control_Array769 <= std_logic_vector(tmp_nfa_dfa_Control_Array(769));
    nfa_dfa_Control_Array770 <= std_logic_vector(tmp_nfa_dfa_Control_Array(770));
    nfa_dfa_Control_Array771 <= std_logic_vector(tmp_nfa_dfa_Control_Array(771));
    nfa_dfa_Control_Array772 <= std_logic_vector(tmp_nfa_dfa_Control_Array(772));
    nfa_dfa_Control_Array773 <= std_logic_vector(tmp_nfa_dfa_Control_Array(773));
    nfa_dfa_Control_Array774 <= std_logic_vector(tmp_nfa_dfa_Control_Array(774));
    nfa_dfa_Control_Array775 <= std_logic_vector(tmp_nfa_dfa_Control_Array(775));
    nfa_dfa_Control_Array776 <= std_logic_vector(tmp_nfa_dfa_Control_Array(776));
    nfa_dfa_Control_Array777 <= std_logic_vector(tmp_nfa_dfa_Control_Array(777));
    nfa_dfa_Control_Array778 <= std_logic_vector(tmp_nfa_dfa_Control_Array(778));
    nfa_dfa_Control_Array779 <= std_logic_vector(tmp_nfa_dfa_Control_Array(779));
    nfa_dfa_Control_Array780 <= std_logic_vector(tmp_nfa_dfa_Control_Array(780));
    nfa_dfa_Control_Array781 <= std_logic_vector(tmp_nfa_dfa_Control_Array(781));
    nfa_dfa_Control_Array782 <= std_logic_vector(tmp_nfa_dfa_Control_Array(782));
    nfa_dfa_Control_Array783 <= std_logic_vector(tmp_nfa_dfa_Control_Array(783));
    nfa_dfa_Control_Array784 <= std_logic_vector(tmp_nfa_dfa_Control_Array(784));
    nfa_dfa_Control_Array785 <= std_logic_vector(tmp_nfa_dfa_Control_Array(785));
    nfa_dfa_Control_Array786 <= std_logic_vector(tmp_nfa_dfa_Control_Array(786));
    nfa_dfa_Control_Array787 <= std_logic_vector(tmp_nfa_dfa_Control_Array(787));
    nfa_dfa_Control_Array788 <= std_logic_vector(tmp_nfa_dfa_Control_Array(788));
    nfa_dfa_Control_Array789 <= std_logic_vector(tmp_nfa_dfa_Control_Array(789));
    nfa_dfa_Control_Array790 <= std_logic_vector(tmp_nfa_dfa_Control_Array(790));
    nfa_dfa_Control_Array791 <= std_logic_vector(tmp_nfa_dfa_Control_Array(791));
    nfa_dfa_Control_Array792 <= std_logic_vector(tmp_nfa_dfa_Control_Array(792));
    nfa_dfa_Control_Array793 <= std_logic_vector(tmp_nfa_dfa_Control_Array(793));
    nfa_dfa_Control_Array794 <= std_logic_vector(tmp_nfa_dfa_Control_Array(794));
    nfa_dfa_Control_Array795 <= std_logic_vector(tmp_nfa_dfa_Control_Array(795));
    nfa_dfa_Control_Array796 <= std_logic_vector(tmp_nfa_dfa_Control_Array(796));
    nfa_dfa_Control_Array797 <= std_logic_vector(tmp_nfa_dfa_Control_Array(797));
    nfa_dfa_Control_Array798 <= std_logic_vector(tmp_nfa_dfa_Control_Array(798));
    nfa_dfa_Control_Array799 <= std_logic_vector(tmp_nfa_dfa_Control_Array(799));
    nfa_dfa_Control_Array800 <= std_logic_vector(tmp_nfa_dfa_Control_Array(800));
    nfa_dfa_Control_Array801 <= std_logic_vector(tmp_nfa_dfa_Control_Array(801));
    nfa_dfa_Control_Array802 <= std_logic_vector(tmp_nfa_dfa_Control_Array(802));
    nfa_dfa_Control_Array803 <= std_logic_vector(tmp_nfa_dfa_Control_Array(803));
    nfa_dfa_Control_Array804 <= std_logic_vector(tmp_nfa_dfa_Control_Array(804));
    nfa_dfa_Control_Array805 <= std_logic_vector(tmp_nfa_dfa_Control_Array(805));
    nfa_dfa_Control_Array806 <= std_logic_vector(tmp_nfa_dfa_Control_Array(806));
    nfa_dfa_Control_Array807 <= std_logic_vector(tmp_nfa_dfa_Control_Array(807));
    nfa_dfa_Control_Array808 <= std_logic_vector(tmp_nfa_dfa_Control_Array(808));
    nfa_dfa_Control_Array809 <= std_logic_vector(tmp_nfa_dfa_Control_Array(809));
    nfa_dfa_Control_Array810 <= std_logic_vector(tmp_nfa_dfa_Control_Array(810));
    nfa_dfa_Control_Array811 <= std_logic_vector(tmp_nfa_dfa_Control_Array(811));
    nfa_dfa_Control_Array812 <= std_logic_vector(tmp_nfa_dfa_Control_Array(812));
    nfa_dfa_Control_Array813 <= std_logic_vector(tmp_nfa_dfa_Control_Array(813));
    nfa_dfa_Control_Array814 <= std_logic_vector(tmp_nfa_dfa_Control_Array(814));
    nfa_dfa_Control_Array815 <= std_logic_vector(tmp_nfa_dfa_Control_Array(815));
    nfa_dfa_Control_Array816 <= std_logic_vector(tmp_nfa_dfa_Control_Array(816));
    nfa_dfa_Control_Array817 <= std_logic_vector(tmp_nfa_dfa_Control_Array(817));
    nfa_dfa_Control_Array818 <= std_logic_vector(tmp_nfa_dfa_Control_Array(818));
    nfa_dfa_Control_Array819 <= std_logic_vector(tmp_nfa_dfa_Control_Array(819));
    nfa_dfa_Control_Array820 <= std_logic_vector(tmp_nfa_dfa_Control_Array(820));
    nfa_dfa_Control_Array821 <= std_logic_vector(tmp_nfa_dfa_Control_Array(821));
    nfa_dfa_Control_Array822 <= std_logic_vector(tmp_nfa_dfa_Control_Array(822));
    nfa_dfa_Control_Array823 <= std_logic_vector(tmp_nfa_dfa_Control_Array(823));
    nfa_dfa_Control_Array824 <= std_logic_vector(tmp_nfa_dfa_Control_Array(824));
    nfa_dfa_Control_Array825 <= std_logic_vector(tmp_nfa_dfa_Control_Array(825));
    nfa_dfa_Control_Array826 <= std_logic_vector(tmp_nfa_dfa_Control_Array(826));
    nfa_dfa_Control_Array827 <= std_logic_vector(tmp_nfa_dfa_Control_Array(827));
    nfa_dfa_Control_Array828 <= std_logic_vector(tmp_nfa_dfa_Control_Array(828));
    nfa_dfa_Control_Array829 <= std_logic_vector(tmp_nfa_dfa_Control_Array(829));
    nfa_dfa_Control_Array830 <= std_logic_vector(tmp_nfa_dfa_Control_Array(830));
    nfa_dfa_Control_Array831 <= std_logic_vector(tmp_nfa_dfa_Control_Array(831));
    nfa_dfa_Control_Array832 <= std_logic_vector(tmp_nfa_dfa_Control_Array(832));
    nfa_dfa_Control_Array833 <= std_logic_vector(tmp_nfa_dfa_Control_Array(833));
    nfa_dfa_Control_Array834 <= std_logic_vector(tmp_nfa_dfa_Control_Array(834));
    nfa_dfa_Control_Array835 <= std_logic_vector(tmp_nfa_dfa_Control_Array(835));
    nfa_dfa_Control_Array836 <= std_logic_vector(tmp_nfa_dfa_Control_Array(836));
    nfa_dfa_Control_Array837 <= std_logic_vector(tmp_nfa_dfa_Control_Array(837));
    nfa_dfa_Control_Array838 <= std_logic_vector(tmp_nfa_dfa_Control_Array(838));
    nfa_dfa_Control_Array839 <= std_logic_vector(tmp_nfa_dfa_Control_Array(839));
    nfa_dfa_Control_Array840 <= std_logic_vector(tmp_nfa_dfa_Control_Array(840));
    nfa_dfa_Control_Array841 <= std_logic_vector(tmp_nfa_dfa_Control_Array(841));
    nfa_dfa_Control_Array842 <= std_logic_vector(tmp_nfa_dfa_Control_Array(842));
    nfa_dfa_Control_Array843 <= std_logic_vector(tmp_nfa_dfa_Control_Array(843));
    nfa_dfa_Control_Array844 <= std_logic_vector(tmp_nfa_dfa_Control_Array(844));
    nfa_dfa_Control_Array845 <= std_logic_vector(tmp_nfa_dfa_Control_Array(845));
    nfa_dfa_Control_Array846 <= std_logic_vector(tmp_nfa_dfa_Control_Array(846));
    nfa_dfa_Control_Array847 <= std_logic_vector(tmp_nfa_dfa_Control_Array(847));
    nfa_dfa_Control_Array848 <= std_logic_vector(tmp_nfa_dfa_Control_Array(848));
    nfa_dfa_Control_Array849 <= std_logic_vector(tmp_nfa_dfa_Control_Array(849));
    nfa_dfa_Control_Array850 <= std_logic_vector(tmp_nfa_dfa_Control_Array(850));
    nfa_dfa_Control_Array851 <= std_logic_vector(tmp_nfa_dfa_Control_Array(851));
    nfa_dfa_Control_Array852 <= std_logic_vector(tmp_nfa_dfa_Control_Array(852));
    nfa_dfa_Control_Array853 <= std_logic_vector(tmp_nfa_dfa_Control_Array(853));
    nfa_dfa_Control_Array854 <= std_logic_vector(tmp_nfa_dfa_Control_Array(854));
    nfa_dfa_Control_Array855 <= std_logic_vector(tmp_nfa_dfa_Control_Array(855));
    nfa_dfa_Control_Array856 <= std_logic_vector(tmp_nfa_dfa_Control_Array(856));
    nfa_dfa_Control_Array857 <= std_logic_vector(tmp_nfa_dfa_Control_Array(857));
    nfa_dfa_Control_Array858 <= std_logic_vector(tmp_nfa_dfa_Control_Array(858));
    nfa_dfa_Control_Array859 <= std_logic_vector(tmp_nfa_dfa_Control_Array(859));
    nfa_dfa_Control_Array860 <= std_logic_vector(tmp_nfa_dfa_Control_Array(860));
    nfa_dfa_Control_Array861 <= std_logic_vector(tmp_nfa_dfa_Control_Array(861));
    nfa_dfa_Control_Array862 <= std_logic_vector(tmp_nfa_dfa_Control_Array(862));
    nfa_dfa_Control_Array863 <= std_logic_vector(tmp_nfa_dfa_Control_Array(863));
    nfa_dfa_Control_Array864 <= std_logic_vector(tmp_nfa_dfa_Control_Array(864));
    nfa_dfa_Control_Array865 <= std_logic_vector(tmp_nfa_dfa_Control_Array(865));
    nfa_dfa_Control_Array866 <= std_logic_vector(tmp_nfa_dfa_Control_Array(866));
    nfa_dfa_Control_Array867 <= std_logic_vector(tmp_nfa_dfa_Control_Array(867));
    nfa_dfa_Control_Array868 <= std_logic_vector(tmp_nfa_dfa_Control_Array(868));
    nfa_dfa_Control_Array869 <= std_logic_vector(tmp_nfa_dfa_Control_Array(869));
    nfa_dfa_Control_Array870 <= std_logic_vector(tmp_nfa_dfa_Control_Array(870));
    nfa_dfa_Control_Array871 <= std_logic_vector(tmp_nfa_dfa_Control_Array(871));
    nfa_dfa_Control_Array872 <= std_logic_vector(tmp_nfa_dfa_Control_Array(872));
    nfa_dfa_Control_Array873 <= std_logic_vector(tmp_nfa_dfa_Control_Array(873));
    nfa_dfa_Control_Array874 <= std_logic_vector(tmp_nfa_dfa_Control_Array(874));
    nfa_dfa_Control_Array875 <= std_logic_vector(tmp_nfa_dfa_Control_Array(875));
    nfa_dfa_Control_Array876 <= std_logic_vector(tmp_nfa_dfa_Control_Array(876));
    nfa_dfa_Control_Array877 <= std_logic_vector(tmp_nfa_dfa_Control_Array(877));
    nfa_dfa_Control_Array878 <= std_logic_vector(tmp_nfa_dfa_Control_Array(878));
    nfa_dfa_Control_Array879 <= std_logic_vector(tmp_nfa_dfa_Control_Array(879));
    nfa_dfa_Control_Array880 <= std_logic_vector(tmp_nfa_dfa_Control_Array(880));
    nfa_dfa_Control_Array881 <= std_logic_vector(tmp_nfa_dfa_Control_Array(881));
    nfa_dfa_Control_Array882 <= std_logic_vector(tmp_nfa_dfa_Control_Array(882));
    nfa_dfa_Control_Array883 <= std_logic_vector(tmp_nfa_dfa_Control_Array(883));
    nfa_dfa_Control_Array884 <= std_logic_vector(tmp_nfa_dfa_Control_Array(884));
    nfa_dfa_Control_Array885 <= std_logic_vector(tmp_nfa_dfa_Control_Array(885));
    nfa_dfa_Control_Array886 <= std_logic_vector(tmp_nfa_dfa_Control_Array(886));
    nfa_dfa_Control_Array887 <= std_logic_vector(tmp_nfa_dfa_Control_Array(887));
    nfa_dfa_Control_Array888 <= std_logic_vector(tmp_nfa_dfa_Control_Array(888));
    nfa_dfa_Control_Array889 <= std_logic_vector(tmp_nfa_dfa_Control_Array(889));
    nfa_dfa_Control_Array890 <= std_logic_vector(tmp_nfa_dfa_Control_Array(890));
    nfa_dfa_Control_Array891 <= std_logic_vector(tmp_nfa_dfa_Control_Array(891));
    nfa_dfa_Control_Array892 <= std_logic_vector(tmp_nfa_dfa_Control_Array(892));
    nfa_dfa_Control_Array893 <= std_logic_vector(tmp_nfa_dfa_Control_Array(893));
    nfa_dfa_Control_Array894 <= std_logic_vector(tmp_nfa_dfa_Control_Array(894));
    nfa_dfa_Control_Array895 <= std_logic_vector(tmp_nfa_dfa_Control_Array(895));
    nfa_dfa_Control_Array896 <= std_logic_vector(tmp_nfa_dfa_Control_Array(896));
    nfa_dfa_Control_Array897 <= std_logic_vector(tmp_nfa_dfa_Control_Array(897));
    nfa_dfa_Control_Array898 <= std_logic_vector(tmp_nfa_dfa_Control_Array(898));
    nfa_dfa_Control_Array899 <= std_logic_vector(tmp_nfa_dfa_Control_Array(899));
    nfa_dfa_Control_Array900 <= std_logic_vector(tmp_nfa_dfa_Control_Array(900));
    nfa_dfa_Control_Array901 <= std_logic_vector(tmp_nfa_dfa_Control_Array(901));
    nfa_dfa_Control_Array902 <= std_logic_vector(tmp_nfa_dfa_Control_Array(902));
    nfa_dfa_Control_Array903 <= std_logic_vector(tmp_nfa_dfa_Control_Array(903));
    nfa_dfa_Control_Array904 <= std_logic_vector(tmp_nfa_dfa_Control_Array(904));
    nfa_dfa_Control_Array905 <= std_logic_vector(tmp_nfa_dfa_Control_Array(905));
    nfa_dfa_Control_Array906 <= std_logic_vector(tmp_nfa_dfa_Control_Array(906));
    nfa_dfa_Control_Array907 <= std_logic_vector(tmp_nfa_dfa_Control_Array(907));
    nfa_dfa_Control_Array908 <= std_logic_vector(tmp_nfa_dfa_Control_Array(908));
    nfa_dfa_Control_Array909 <= std_logic_vector(tmp_nfa_dfa_Control_Array(909));
    nfa_dfa_Control_Array910 <= std_logic_vector(tmp_nfa_dfa_Control_Array(910));
    nfa_dfa_Control_Array911 <= std_logic_vector(tmp_nfa_dfa_Control_Array(911));
    nfa_dfa_Control_Array912 <= std_logic_vector(tmp_nfa_dfa_Control_Array(912));
    nfa_dfa_Control_Array913 <= std_logic_vector(tmp_nfa_dfa_Control_Array(913));
    nfa_dfa_Control_Array914 <= std_logic_vector(tmp_nfa_dfa_Control_Array(914));
    nfa_dfa_Control_Array915 <= std_logic_vector(tmp_nfa_dfa_Control_Array(915));
    nfa_dfa_Control_Array916 <= std_logic_vector(tmp_nfa_dfa_Control_Array(916));
    nfa_dfa_Control_Array917 <= std_logic_vector(tmp_nfa_dfa_Control_Array(917));
    nfa_dfa_Control_Array918 <= std_logic_vector(tmp_nfa_dfa_Control_Array(918));
    nfa_dfa_Control_Array919 <= std_logic_vector(tmp_nfa_dfa_Control_Array(919));
    nfa_dfa_Control_Array920 <= std_logic_vector(tmp_nfa_dfa_Control_Array(920));
    nfa_dfa_Control_Array921 <= std_logic_vector(tmp_nfa_dfa_Control_Array(921));
    nfa_dfa_Control_Array922 <= std_logic_vector(tmp_nfa_dfa_Control_Array(922));
    nfa_dfa_Control_Array923 <= std_logic_vector(tmp_nfa_dfa_Control_Array(923));
    nfa_dfa_Control_Array924 <= std_logic_vector(tmp_nfa_dfa_Control_Array(924));
    nfa_dfa_Control_Array925 <= std_logic_vector(tmp_nfa_dfa_Control_Array(925));
    nfa_dfa_Control_Array926 <= std_logic_vector(tmp_nfa_dfa_Control_Array(926));
    nfa_dfa_Control_Array927 <= std_logic_vector(tmp_nfa_dfa_Control_Array(927));
    nfa_dfa_Control_Array928 <= std_logic_vector(tmp_nfa_dfa_Control_Array(928));
    nfa_dfa_Control_Array929 <= std_logic_vector(tmp_nfa_dfa_Control_Array(929));
    nfa_dfa_Control_Array930 <= std_logic_vector(tmp_nfa_dfa_Control_Array(930));
    nfa_dfa_Control_Array931 <= std_logic_vector(tmp_nfa_dfa_Control_Array(931));
    nfa_dfa_Control_Array932 <= std_logic_vector(tmp_nfa_dfa_Control_Array(932));
    nfa_dfa_Control_Array933 <= std_logic_vector(tmp_nfa_dfa_Control_Array(933));
    nfa_dfa_Control_Array934 <= std_logic_vector(tmp_nfa_dfa_Control_Array(934));
    nfa_dfa_Control_Array935 <= std_logic_vector(tmp_nfa_dfa_Control_Array(935));
    nfa_dfa_Control_Array936 <= std_logic_vector(tmp_nfa_dfa_Control_Array(936));
    nfa_dfa_Control_Array937 <= std_logic_vector(tmp_nfa_dfa_Control_Array(937));
    nfa_dfa_Control_Array938 <= std_logic_vector(tmp_nfa_dfa_Control_Array(938));
    nfa_dfa_Control_Array939 <= std_logic_vector(tmp_nfa_dfa_Control_Array(939));
    nfa_dfa_Control_Array940 <= std_logic_vector(tmp_nfa_dfa_Control_Array(940));
    nfa_dfa_Control_Array941 <= std_logic_vector(tmp_nfa_dfa_Control_Array(941));
    nfa_dfa_Control_Array942 <= std_logic_vector(tmp_nfa_dfa_Control_Array(942));
    nfa_dfa_Control_Array943 <= std_logic_vector(tmp_nfa_dfa_Control_Array(943));
    nfa_dfa_Control_Array944 <= std_logic_vector(tmp_nfa_dfa_Control_Array(944));
    nfa_dfa_Control_Array945 <= std_logic_vector(tmp_nfa_dfa_Control_Array(945));
    nfa_dfa_Control_Array946 <= std_logic_vector(tmp_nfa_dfa_Control_Array(946));
    nfa_dfa_Control_Array947 <= std_logic_vector(tmp_nfa_dfa_Control_Array(947));
    nfa_dfa_Control_Array948 <= std_logic_vector(tmp_nfa_dfa_Control_Array(948));
    nfa_dfa_Control_Array949 <= std_logic_vector(tmp_nfa_dfa_Control_Array(949));
    nfa_dfa_Control_Array950 <= std_logic_vector(tmp_nfa_dfa_Control_Array(950));
    nfa_dfa_Control_Array951 <= std_logic_vector(tmp_nfa_dfa_Control_Array(951));
    nfa_dfa_Control_Array952 <= std_logic_vector(tmp_nfa_dfa_Control_Array(952));
    nfa_dfa_Control_Array953 <= std_logic_vector(tmp_nfa_dfa_Control_Array(953));
    nfa_dfa_Control_Array954 <= std_logic_vector(tmp_nfa_dfa_Control_Array(954));
    nfa_dfa_Control_Array955 <= std_logic_vector(tmp_nfa_dfa_Control_Array(955));
    nfa_dfa_Control_Array956 <= std_logic_vector(tmp_nfa_dfa_Control_Array(956));
    nfa_dfa_Control_Array957 <= std_logic_vector(tmp_nfa_dfa_Control_Array(957));
    nfa_dfa_Control_Array958 <= std_logic_vector(tmp_nfa_dfa_Control_Array(958));
    nfa_dfa_Control_Array959 <= std_logic_vector(tmp_nfa_dfa_Control_Array(959));
    nfa_dfa_Control_Array960 <= std_logic_vector(tmp_nfa_dfa_Control_Array(960));
    nfa_dfa_Control_Array961 <= std_logic_vector(tmp_nfa_dfa_Control_Array(961));
    nfa_dfa_Control_Array962 <= std_logic_vector(tmp_nfa_dfa_Control_Array(962));
    nfa_dfa_Control_Array963 <= std_logic_vector(tmp_nfa_dfa_Control_Array(963));
    nfa_dfa_Control_Array964 <= std_logic_vector(tmp_nfa_dfa_Control_Array(964));
    nfa_dfa_Control_Array965 <= std_logic_vector(tmp_nfa_dfa_Control_Array(965));
    nfa_dfa_Control_Array966 <= std_logic_vector(tmp_nfa_dfa_Control_Array(966));
    nfa_dfa_Control_Array967 <= std_logic_vector(tmp_nfa_dfa_Control_Array(967));
    nfa_dfa_Control_Array968 <= std_logic_vector(tmp_nfa_dfa_Control_Array(968));
    nfa_dfa_Control_Array969 <= std_logic_vector(tmp_nfa_dfa_Control_Array(969));
    nfa_dfa_Control_Array970 <= std_logic_vector(tmp_nfa_dfa_Control_Array(970));
    nfa_dfa_Control_Array971 <= std_logic_vector(tmp_nfa_dfa_Control_Array(971));
    nfa_dfa_Control_Array972 <= std_logic_vector(tmp_nfa_dfa_Control_Array(972));
    nfa_dfa_Control_Array973 <= std_logic_vector(tmp_nfa_dfa_Control_Array(973));
    nfa_dfa_Control_Array974 <= std_logic_vector(tmp_nfa_dfa_Control_Array(974));
    nfa_dfa_Control_Array975 <= std_logic_vector(tmp_nfa_dfa_Control_Array(975));
    nfa_dfa_Control_Array976 <= std_logic_vector(tmp_nfa_dfa_Control_Array(976));
    nfa_dfa_Control_Array977 <= std_logic_vector(tmp_nfa_dfa_Control_Array(977));
    nfa_dfa_Control_Array978 <= std_logic_vector(tmp_nfa_dfa_Control_Array(978));
    nfa_dfa_Control_Array979 <= std_logic_vector(tmp_nfa_dfa_Control_Array(979));
    nfa_dfa_Control_Array980 <= std_logic_vector(tmp_nfa_dfa_Control_Array(980));
    nfa_dfa_Control_Array981 <= std_logic_vector(tmp_nfa_dfa_Control_Array(981));
    nfa_dfa_Control_Array982 <= std_logic_vector(tmp_nfa_dfa_Control_Array(982));
    nfa_dfa_Control_Array983 <= std_logic_vector(tmp_nfa_dfa_Control_Array(983));
    nfa_dfa_Control_Array984 <= std_logic_vector(tmp_nfa_dfa_Control_Array(984));
    nfa_dfa_Control_Array985 <= std_logic_vector(tmp_nfa_dfa_Control_Array(985));
    nfa_dfa_Control_Array986 <= std_logic_vector(tmp_nfa_dfa_Control_Array(986));
    nfa_dfa_Control_Array987 <= std_logic_vector(tmp_nfa_dfa_Control_Array(987));
    nfa_dfa_Control_Array988 <= std_logic_vector(tmp_nfa_dfa_Control_Array(988));
    nfa_dfa_Control_Array989 <= std_logic_vector(tmp_nfa_dfa_Control_Array(989));
    nfa_dfa_Control_Array990 <= std_logic_vector(tmp_nfa_dfa_Control_Array(990));
    nfa_dfa_Control_Array991 <= std_logic_vector(tmp_nfa_dfa_Control_Array(991));
    nfa_dfa_Control_Array992 <= std_logic_vector(tmp_nfa_dfa_Control_Array(992));
    nfa_dfa_Control_Array993 <= std_logic_vector(tmp_nfa_dfa_Control_Array(993));
    nfa_dfa_Control_Array994 <= std_logic_vector(tmp_nfa_dfa_Control_Array(994));
    nfa_dfa_Control_Array995 <= std_logic_vector(tmp_nfa_dfa_Control_Array(995));
    nfa_dfa_Control_Array996 <= std_logic_vector(tmp_nfa_dfa_Control_Array(996));
    nfa_dfa_Control_Array997 <= std_logic_vector(tmp_nfa_dfa_Control_Array(997));
    nfa_dfa_Control_Array998 <= std_logic_vector(tmp_nfa_dfa_Control_Array(998));
    nfa_dfa_Control_Array999 <= std_logic_vector(tmp_nfa_dfa_Control_Array(999));

    -- Entity sme_intro signals
    sme_intro: entity work.sme_intro
    port map (
        -- Output bus nfa_dfa_Control
        nfa_dfa_Control_Valid => nfa_dfa_Control_Valid,
        nfa_dfa_Control_Reset => nfa_dfa_Control_Reset,
        nfa_dfa_Control_Length => tmp_nfa_dfa_Control_Length,
        nfa_dfa_Control_Array => tmp_nfa_dfa_Control_Array,

        -- Input bus nfa_dfa_Traversal
        nfa_dfa_Traversal_Valid => nfa_dfa_Traversal_Valid,

        ENB => ENB,
        RST => RST,
        FIN => FIN,
        CLK => CLK
    );

-- User defined processes here
-- #### USER-DATA-CODE-START
-- #### USER-DATA-CODE-END

end RTL;