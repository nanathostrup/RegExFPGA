library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- library SYSTEM_TYPES;
use work.SYSTEM_TYPES.ALL;

-- library CUSTOM_TYPES;
use work.CUSTOM_TYPES.ALL;

-- User defined packages here
-- #### USER-DATA-IMPORTS-START
-- #### USER-DATA-IMPORTS-END

entity sme_intro_export is
    port(
        -- Top-level bus Control signals
        Control_Valid: out STD_LOGIC;
        Control_Reset: out STD_LOGIC;
        Control_Length: out STD_LOGIC_VECTOR(31 downto 0);
        Control_Array0: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array1: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array2: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array3: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array4: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array5: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array6: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array7: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array8: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array9: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array10: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array11: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array12: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array13: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array14: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array15: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array16: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array17: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array18: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array19: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array20: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array21: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array22: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array23: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array24: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array25: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array26: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array27: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array28: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array29: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array30: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array31: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array32: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array33: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array34: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array35: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array36: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array37: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array38: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array39: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array40: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array41: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array42: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array43: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array44: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array45: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array46: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array47: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array48: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array49: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array50: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array51: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array52: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array53: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array54: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array55: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array56: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array57: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array58: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array59: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array60: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array61: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array62: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array63: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array64: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array65: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array66: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array67: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array68: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array69: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array70: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array71: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array72: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array73: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array74: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array75: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array76: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array77: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array78: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array79: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array80: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array81: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array82: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array83: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array84: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array85: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array86: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array87: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array88: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array89: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array90: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array91: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array92: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array93: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array94: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array95: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array96: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array97: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array98: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array99: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array100: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array101: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array102: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array103: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array104: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array105: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array106: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array107: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array108: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array109: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array110: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array111: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array112: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array113: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array114: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array115: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array116: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array117: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array118: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array119: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array120: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array121: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array122: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array123: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array124: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array125: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array126: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array127: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array128: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array129: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array130: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array131: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array132: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array133: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array134: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array135: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array136: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array137: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array138: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array139: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array140: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array141: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array142: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array143: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array144: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array145: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array146: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array147: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array148: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array149: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array150: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array151: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array152: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array153: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array154: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array155: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array156: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array157: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array158: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array159: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array160: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array161: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array162: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array163: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array164: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array165: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array166: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array167: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array168: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array169: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array170: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array171: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array172: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array173: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array174: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array175: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array176: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array177: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array178: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array179: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array180: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array181: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array182: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array183: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array184: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array185: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array186: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array187: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array188: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array189: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array190: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array191: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array192: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array193: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array194: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array195: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array196: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array197: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array198: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array199: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array200: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array201: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array202: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array203: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array204: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array205: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array206: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array207: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array208: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array209: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array210: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array211: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array212: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array213: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array214: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array215: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array216: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array217: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array218: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array219: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array220: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array221: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array222: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array223: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array224: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array225: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array226: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array227: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array228: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array229: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array230: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array231: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array232: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array233: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array234: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array235: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array236: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array237: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array238: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array239: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array240: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array241: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array242: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array243: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array244: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array245: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array246: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array247: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array248: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array249: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array250: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array251: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array252: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array253: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array254: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array255: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array256: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array257: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array258: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array259: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array260: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array261: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array262: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array263: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array264: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array265: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array266: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array267: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array268: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array269: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array270: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array271: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array272: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array273: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array274: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array275: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array276: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array277: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array278: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array279: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array280: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array281: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array282: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array283: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array284: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array285: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array286: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array287: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array288: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array289: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array290: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array291: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array292: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array293: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array294: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array295: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array296: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array297: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array298: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array299: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array300: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array301: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array302: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array303: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array304: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array305: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array306: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array307: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array308: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array309: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array310: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array311: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array312: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array313: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array314: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array315: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array316: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array317: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array318: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array319: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array320: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array321: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array322: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array323: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array324: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array325: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array326: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array327: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array328: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array329: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array330: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array331: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array332: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array333: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array334: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array335: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array336: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array337: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array338: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array339: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array340: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array341: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array342: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array343: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array344: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array345: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array346: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array347: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array348: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array349: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array350: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array351: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array352: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array353: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array354: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array355: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array356: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array357: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array358: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array359: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array360: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array361: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array362: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array363: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array364: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array365: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array366: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array367: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array368: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array369: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array370: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array371: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array372: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array373: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array374: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array375: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array376: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array377: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array378: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array379: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array380: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array381: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array382: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array383: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array384: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array385: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array386: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array387: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array388: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array389: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array390: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array391: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array392: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array393: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array394: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array395: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array396: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array397: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array398: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array399: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array400: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array401: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array402: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array403: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array404: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array405: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array406: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array407: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array408: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array409: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array410: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array411: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array412: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array413: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array414: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array415: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array416: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array417: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array418: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array419: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array420: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array421: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array422: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array423: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array424: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array425: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array426: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array427: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array428: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array429: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array430: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array431: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array432: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array433: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array434: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array435: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array436: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array437: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array438: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array439: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array440: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array441: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array442: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array443: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array444: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array445: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array446: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array447: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array448: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array449: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array450: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array451: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array452: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array453: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array454: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array455: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array456: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array457: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array458: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array459: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array460: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array461: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array462: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array463: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array464: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array465: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array466: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array467: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array468: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array469: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array470: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array471: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array472: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array473: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array474: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array475: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array476: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array477: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array478: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array479: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array480: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array481: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array482: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array483: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array484: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array485: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array486: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array487: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array488: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array489: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array490: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array491: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array492: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array493: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array494: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array495: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array496: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array497: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array498: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array499: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array500: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array501: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array502: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array503: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array504: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array505: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array506: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array507: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array508: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array509: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array510: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array511: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array512: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array513: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array514: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array515: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array516: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array517: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array518: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array519: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array520: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array521: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array522: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array523: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array524: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array525: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array526: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array527: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array528: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array529: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array530: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array531: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array532: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array533: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array534: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array535: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array536: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array537: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array538: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array539: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array540: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array541: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array542: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array543: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array544: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array545: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array546: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array547: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array548: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array549: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array550: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array551: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array552: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array553: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array554: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array555: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array556: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array557: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array558: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array559: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array560: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array561: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array562: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array563: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array564: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array565: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array566: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array567: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array568: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array569: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array570: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array571: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array572: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array573: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array574: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array575: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array576: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array577: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array578: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array579: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array580: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array581: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array582: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array583: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array584: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array585: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array586: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array587: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array588: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array589: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array590: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array591: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array592: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array593: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array594: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array595: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array596: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array597: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array598: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array599: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array600: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array601: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array602: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array603: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array604: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array605: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array606: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array607: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array608: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array609: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array610: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array611: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array612: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array613: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array614: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array615: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array616: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array617: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array618: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array619: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array620: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array621: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array622: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array623: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array624: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array625: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array626: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array627: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array628: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array629: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array630: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array631: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array632: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array633: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array634: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array635: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array636: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array637: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array638: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array639: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array640: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array641: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array642: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array643: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array644: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array645: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array646: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array647: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array648: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array649: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array650: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array651: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array652: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array653: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array654: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array655: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array656: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array657: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array658: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array659: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array660: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array661: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array662: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array663: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array664: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array665: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array666: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array667: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array668: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array669: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array670: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array671: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array672: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array673: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array674: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array675: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array676: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array677: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array678: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array679: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array680: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array681: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array682: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array683: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array684: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array685: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array686: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array687: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array688: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array689: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array690: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array691: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array692: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array693: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array694: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array695: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array696: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array697: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array698: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array699: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array700: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array701: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array702: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array703: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array704: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array705: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array706: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array707: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array708: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array709: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array710: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array711: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array712: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array713: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array714: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array715: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array716: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array717: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array718: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array719: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array720: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array721: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array722: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array723: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array724: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array725: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array726: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array727: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array728: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array729: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array730: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array731: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array732: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array733: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array734: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array735: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array736: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array737: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array738: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array739: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array740: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array741: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array742: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array743: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array744: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array745: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array746: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array747: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array748: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array749: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array750: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array751: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array752: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array753: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array754: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array755: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array756: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array757: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array758: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array759: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array760: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array761: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array762: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array763: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array764: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array765: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array766: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array767: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array768: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array769: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array770: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array771: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array772: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array773: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array774: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array775: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array776: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array777: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array778: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array779: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array780: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array781: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array782: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array783: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array784: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array785: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array786: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array787: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array788: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array789: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array790: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array791: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array792: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array793: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array794: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array795: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array796: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array797: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array798: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array799: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array800: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array801: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array802: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array803: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array804: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array805: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array806: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array807: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array808: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array809: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array810: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array811: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array812: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array813: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array814: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array815: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array816: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array817: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array818: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array819: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array820: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array821: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array822: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array823: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array824: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array825: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array826: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array827: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array828: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array829: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array830: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array831: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array832: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array833: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array834: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array835: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array836: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array837: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array838: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array839: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array840: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array841: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array842: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array843: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array844: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array845: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array846: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array847: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array848: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array849: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array850: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array851: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array852: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array853: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array854: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array855: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array856: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array857: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array858: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array859: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array860: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array861: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array862: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array863: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array864: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array865: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array866: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array867: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array868: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array869: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array870: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array871: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array872: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array873: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array874: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array875: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array876: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array877: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array878: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array879: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array880: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array881: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array882: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array883: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array884: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array885: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array886: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array887: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array888: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array889: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array890: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array891: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array892: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array893: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array894: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array895: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array896: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array897: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array898: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array899: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array900: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array901: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array902: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array903: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array904: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array905: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array906: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array907: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array908: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array909: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array910: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array911: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array912: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array913: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array914: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array915: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array916: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array917: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array918: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array919: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array920: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array921: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array922: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array923: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array924: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array925: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array926: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array927: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array928: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array929: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array930: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array931: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array932: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array933: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array934: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array935: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array936: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array937: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array938: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array939: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array940: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array941: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array942: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array943: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array944: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array945: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array946: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array947: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array948: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array949: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array950: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array951: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array952: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array953: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array954: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array955: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array956: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array957: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array958: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array959: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array960: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array961: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array962: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array963: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array964: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array965: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array966: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array967: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array968: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array969: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array970: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array971: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array972: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array973: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array974: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array975: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array976: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array977: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array978: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array979: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array980: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array981: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array982: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array983: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array984: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array985: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array986: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array987: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array988: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array989: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array990: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array991: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array992: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array993: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array994: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array995: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array996: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array997: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array998: out STD_LOGIC_VECTOR(7 downto 0);
        Control_Array999: out STD_LOGIC_VECTOR(7 downto 0);

        -- Top-level bus Traversal signals
        Traversal_Valid: in STD_LOGIC;

        -- User defined signals here
        -- #### USER-DATA-ENTITYSIGNALS-START
        -- #### USER-DATA-ENTITYSIGNALS-END

        -- Enable signal
        ENB : in STD_LOGIC;

        -- Reset signal
        RST : in STD_LOGIC;

        -- Finished signal
        FIN : out Std_logic;

        -- Clock signal
        CLK : in STD_LOGIC
    );
end sme_intro_export;

architecture RTL of sme_intro_export is

    -- User defined signals here
    -- #### USER-DATA-SIGNALS-START
    -- #### USER-DATA-SIGNALS-END

    -- Intermediate conversion signal to convert internal types to external ones
    signal tmp_Control_Length : T_SYSTEM_INT32;
    signal tmp_Control_Array : Control_Array_type;

begin

    -- Carry converted signals from entity to wrapped outputs
    Control_Length <= std_logic_vector(tmp_Control_Length);
    Control_Array0 <= std_logic_vector(tmp_Control_Array(0));
    Control_Array1 <= std_logic_vector(tmp_Control_Array(1));
    Control_Array2 <= std_logic_vector(tmp_Control_Array(2));
    Control_Array3 <= std_logic_vector(tmp_Control_Array(3));
    Control_Array4 <= std_logic_vector(tmp_Control_Array(4));
    Control_Array5 <= std_logic_vector(tmp_Control_Array(5));
    Control_Array6 <= std_logic_vector(tmp_Control_Array(6));
    Control_Array7 <= std_logic_vector(tmp_Control_Array(7));
    Control_Array8 <= std_logic_vector(tmp_Control_Array(8));
    Control_Array9 <= std_logic_vector(tmp_Control_Array(9));
    Control_Array10 <= std_logic_vector(tmp_Control_Array(10));
    Control_Array11 <= std_logic_vector(tmp_Control_Array(11));
    Control_Array12 <= std_logic_vector(tmp_Control_Array(12));
    Control_Array13 <= std_logic_vector(tmp_Control_Array(13));
    Control_Array14 <= std_logic_vector(tmp_Control_Array(14));
    Control_Array15 <= std_logic_vector(tmp_Control_Array(15));
    Control_Array16 <= std_logic_vector(tmp_Control_Array(16));
    Control_Array17 <= std_logic_vector(tmp_Control_Array(17));
    Control_Array18 <= std_logic_vector(tmp_Control_Array(18));
    Control_Array19 <= std_logic_vector(tmp_Control_Array(19));
    Control_Array20 <= std_logic_vector(tmp_Control_Array(20));
    Control_Array21 <= std_logic_vector(tmp_Control_Array(21));
    Control_Array22 <= std_logic_vector(tmp_Control_Array(22));
    Control_Array23 <= std_logic_vector(tmp_Control_Array(23));
    Control_Array24 <= std_logic_vector(tmp_Control_Array(24));
    Control_Array25 <= std_logic_vector(tmp_Control_Array(25));
    Control_Array26 <= std_logic_vector(tmp_Control_Array(26));
    Control_Array27 <= std_logic_vector(tmp_Control_Array(27));
    Control_Array28 <= std_logic_vector(tmp_Control_Array(28));
    Control_Array29 <= std_logic_vector(tmp_Control_Array(29));
    Control_Array30 <= std_logic_vector(tmp_Control_Array(30));
    Control_Array31 <= std_logic_vector(tmp_Control_Array(31));
    Control_Array32 <= std_logic_vector(tmp_Control_Array(32));
    Control_Array33 <= std_logic_vector(tmp_Control_Array(33));
    Control_Array34 <= std_logic_vector(tmp_Control_Array(34));
    Control_Array35 <= std_logic_vector(tmp_Control_Array(35));
    Control_Array36 <= std_logic_vector(tmp_Control_Array(36));
    Control_Array37 <= std_logic_vector(tmp_Control_Array(37));
    Control_Array38 <= std_logic_vector(tmp_Control_Array(38));
    Control_Array39 <= std_logic_vector(tmp_Control_Array(39));
    Control_Array40 <= std_logic_vector(tmp_Control_Array(40));
    Control_Array41 <= std_logic_vector(tmp_Control_Array(41));
    Control_Array42 <= std_logic_vector(tmp_Control_Array(42));
    Control_Array43 <= std_logic_vector(tmp_Control_Array(43));
    Control_Array44 <= std_logic_vector(tmp_Control_Array(44));
    Control_Array45 <= std_logic_vector(tmp_Control_Array(45));
    Control_Array46 <= std_logic_vector(tmp_Control_Array(46));
    Control_Array47 <= std_logic_vector(tmp_Control_Array(47));
    Control_Array48 <= std_logic_vector(tmp_Control_Array(48));
    Control_Array49 <= std_logic_vector(tmp_Control_Array(49));
    Control_Array50 <= std_logic_vector(tmp_Control_Array(50));
    Control_Array51 <= std_logic_vector(tmp_Control_Array(51));
    Control_Array52 <= std_logic_vector(tmp_Control_Array(52));
    Control_Array53 <= std_logic_vector(tmp_Control_Array(53));
    Control_Array54 <= std_logic_vector(tmp_Control_Array(54));
    Control_Array55 <= std_logic_vector(tmp_Control_Array(55));
    Control_Array56 <= std_logic_vector(tmp_Control_Array(56));
    Control_Array57 <= std_logic_vector(tmp_Control_Array(57));
    Control_Array58 <= std_logic_vector(tmp_Control_Array(58));
    Control_Array59 <= std_logic_vector(tmp_Control_Array(59));
    Control_Array60 <= std_logic_vector(tmp_Control_Array(60));
    Control_Array61 <= std_logic_vector(tmp_Control_Array(61));
    Control_Array62 <= std_logic_vector(tmp_Control_Array(62));
    Control_Array63 <= std_logic_vector(tmp_Control_Array(63));
    Control_Array64 <= std_logic_vector(tmp_Control_Array(64));
    Control_Array65 <= std_logic_vector(tmp_Control_Array(65));
    Control_Array66 <= std_logic_vector(tmp_Control_Array(66));
    Control_Array67 <= std_logic_vector(tmp_Control_Array(67));
    Control_Array68 <= std_logic_vector(tmp_Control_Array(68));
    Control_Array69 <= std_logic_vector(tmp_Control_Array(69));
    Control_Array70 <= std_logic_vector(tmp_Control_Array(70));
    Control_Array71 <= std_logic_vector(tmp_Control_Array(71));
    Control_Array72 <= std_logic_vector(tmp_Control_Array(72));
    Control_Array73 <= std_logic_vector(tmp_Control_Array(73));
    Control_Array74 <= std_logic_vector(tmp_Control_Array(74));
    Control_Array75 <= std_logic_vector(tmp_Control_Array(75));
    Control_Array76 <= std_logic_vector(tmp_Control_Array(76));
    Control_Array77 <= std_logic_vector(tmp_Control_Array(77));
    Control_Array78 <= std_logic_vector(tmp_Control_Array(78));
    Control_Array79 <= std_logic_vector(tmp_Control_Array(79));
    Control_Array80 <= std_logic_vector(tmp_Control_Array(80));
    Control_Array81 <= std_logic_vector(tmp_Control_Array(81));
    Control_Array82 <= std_logic_vector(tmp_Control_Array(82));
    Control_Array83 <= std_logic_vector(tmp_Control_Array(83));
    Control_Array84 <= std_logic_vector(tmp_Control_Array(84));
    Control_Array85 <= std_logic_vector(tmp_Control_Array(85));
    Control_Array86 <= std_logic_vector(tmp_Control_Array(86));
    Control_Array87 <= std_logic_vector(tmp_Control_Array(87));
    Control_Array88 <= std_logic_vector(tmp_Control_Array(88));
    Control_Array89 <= std_logic_vector(tmp_Control_Array(89));
    Control_Array90 <= std_logic_vector(tmp_Control_Array(90));
    Control_Array91 <= std_logic_vector(tmp_Control_Array(91));
    Control_Array92 <= std_logic_vector(tmp_Control_Array(92));
    Control_Array93 <= std_logic_vector(tmp_Control_Array(93));
    Control_Array94 <= std_logic_vector(tmp_Control_Array(94));
    Control_Array95 <= std_logic_vector(tmp_Control_Array(95));
    Control_Array96 <= std_logic_vector(tmp_Control_Array(96));
    Control_Array97 <= std_logic_vector(tmp_Control_Array(97));
    Control_Array98 <= std_logic_vector(tmp_Control_Array(98));
    Control_Array99 <= std_logic_vector(tmp_Control_Array(99));
    Control_Array100 <= std_logic_vector(tmp_Control_Array(100));
    Control_Array101 <= std_logic_vector(tmp_Control_Array(101));
    Control_Array102 <= std_logic_vector(tmp_Control_Array(102));
    Control_Array103 <= std_logic_vector(tmp_Control_Array(103));
    Control_Array104 <= std_logic_vector(tmp_Control_Array(104));
    Control_Array105 <= std_logic_vector(tmp_Control_Array(105));
    Control_Array106 <= std_logic_vector(tmp_Control_Array(106));
    Control_Array107 <= std_logic_vector(tmp_Control_Array(107));
    Control_Array108 <= std_logic_vector(tmp_Control_Array(108));
    Control_Array109 <= std_logic_vector(tmp_Control_Array(109));
    Control_Array110 <= std_logic_vector(tmp_Control_Array(110));
    Control_Array111 <= std_logic_vector(tmp_Control_Array(111));
    Control_Array112 <= std_logic_vector(tmp_Control_Array(112));
    Control_Array113 <= std_logic_vector(tmp_Control_Array(113));
    Control_Array114 <= std_logic_vector(tmp_Control_Array(114));
    Control_Array115 <= std_logic_vector(tmp_Control_Array(115));
    Control_Array116 <= std_logic_vector(tmp_Control_Array(116));
    Control_Array117 <= std_logic_vector(tmp_Control_Array(117));
    Control_Array118 <= std_logic_vector(tmp_Control_Array(118));
    Control_Array119 <= std_logic_vector(tmp_Control_Array(119));
    Control_Array120 <= std_logic_vector(tmp_Control_Array(120));
    Control_Array121 <= std_logic_vector(tmp_Control_Array(121));
    Control_Array122 <= std_logic_vector(tmp_Control_Array(122));
    Control_Array123 <= std_logic_vector(tmp_Control_Array(123));
    Control_Array124 <= std_logic_vector(tmp_Control_Array(124));
    Control_Array125 <= std_logic_vector(tmp_Control_Array(125));
    Control_Array126 <= std_logic_vector(tmp_Control_Array(126));
    Control_Array127 <= std_logic_vector(tmp_Control_Array(127));
    Control_Array128 <= std_logic_vector(tmp_Control_Array(128));
    Control_Array129 <= std_logic_vector(tmp_Control_Array(129));
    Control_Array130 <= std_logic_vector(tmp_Control_Array(130));
    Control_Array131 <= std_logic_vector(tmp_Control_Array(131));
    Control_Array132 <= std_logic_vector(tmp_Control_Array(132));
    Control_Array133 <= std_logic_vector(tmp_Control_Array(133));
    Control_Array134 <= std_logic_vector(tmp_Control_Array(134));
    Control_Array135 <= std_logic_vector(tmp_Control_Array(135));
    Control_Array136 <= std_logic_vector(tmp_Control_Array(136));
    Control_Array137 <= std_logic_vector(tmp_Control_Array(137));
    Control_Array138 <= std_logic_vector(tmp_Control_Array(138));
    Control_Array139 <= std_logic_vector(tmp_Control_Array(139));
    Control_Array140 <= std_logic_vector(tmp_Control_Array(140));
    Control_Array141 <= std_logic_vector(tmp_Control_Array(141));
    Control_Array142 <= std_logic_vector(tmp_Control_Array(142));
    Control_Array143 <= std_logic_vector(tmp_Control_Array(143));
    Control_Array144 <= std_logic_vector(tmp_Control_Array(144));
    Control_Array145 <= std_logic_vector(tmp_Control_Array(145));
    Control_Array146 <= std_logic_vector(tmp_Control_Array(146));
    Control_Array147 <= std_logic_vector(tmp_Control_Array(147));
    Control_Array148 <= std_logic_vector(tmp_Control_Array(148));
    Control_Array149 <= std_logic_vector(tmp_Control_Array(149));
    Control_Array150 <= std_logic_vector(tmp_Control_Array(150));
    Control_Array151 <= std_logic_vector(tmp_Control_Array(151));
    Control_Array152 <= std_logic_vector(tmp_Control_Array(152));
    Control_Array153 <= std_logic_vector(tmp_Control_Array(153));
    Control_Array154 <= std_logic_vector(tmp_Control_Array(154));
    Control_Array155 <= std_logic_vector(tmp_Control_Array(155));
    Control_Array156 <= std_logic_vector(tmp_Control_Array(156));
    Control_Array157 <= std_logic_vector(tmp_Control_Array(157));
    Control_Array158 <= std_logic_vector(tmp_Control_Array(158));
    Control_Array159 <= std_logic_vector(tmp_Control_Array(159));
    Control_Array160 <= std_logic_vector(tmp_Control_Array(160));
    Control_Array161 <= std_logic_vector(tmp_Control_Array(161));
    Control_Array162 <= std_logic_vector(tmp_Control_Array(162));
    Control_Array163 <= std_logic_vector(tmp_Control_Array(163));
    Control_Array164 <= std_logic_vector(tmp_Control_Array(164));
    Control_Array165 <= std_logic_vector(tmp_Control_Array(165));
    Control_Array166 <= std_logic_vector(tmp_Control_Array(166));
    Control_Array167 <= std_logic_vector(tmp_Control_Array(167));
    Control_Array168 <= std_logic_vector(tmp_Control_Array(168));
    Control_Array169 <= std_logic_vector(tmp_Control_Array(169));
    Control_Array170 <= std_logic_vector(tmp_Control_Array(170));
    Control_Array171 <= std_logic_vector(tmp_Control_Array(171));
    Control_Array172 <= std_logic_vector(tmp_Control_Array(172));
    Control_Array173 <= std_logic_vector(tmp_Control_Array(173));
    Control_Array174 <= std_logic_vector(tmp_Control_Array(174));
    Control_Array175 <= std_logic_vector(tmp_Control_Array(175));
    Control_Array176 <= std_logic_vector(tmp_Control_Array(176));
    Control_Array177 <= std_logic_vector(tmp_Control_Array(177));
    Control_Array178 <= std_logic_vector(tmp_Control_Array(178));
    Control_Array179 <= std_logic_vector(tmp_Control_Array(179));
    Control_Array180 <= std_logic_vector(tmp_Control_Array(180));
    Control_Array181 <= std_logic_vector(tmp_Control_Array(181));
    Control_Array182 <= std_logic_vector(tmp_Control_Array(182));
    Control_Array183 <= std_logic_vector(tmp_Control_Array(183));
    Control_Array184 <= std_logic_vector(tmp_Control_Array(184));
    Control_Array185 <= std_logic_vector(tmp_Control_Array(185));
    Control_Array186 <= std_logic_vector(tmp_Control_Array(186));
    Control_Array187 <= std_logic_vector(tmp_Control_Array(187));
    Control_Array188 <= std_logic_vector(tmp_Control_Array(188));
    Control_Array189 <= std_logic_vector(tmp_Control_Array(189));
    Control_Array190 <= std_logic_vector(tmp_Control_Array(190));
    Control_Array191 <= std_logic_vector(tmp_Control_Array(191));
    Control_Array192 <= std_logic_vector(tmp_Control_Array(192));
    Control_Array193 <= std_logic_vector(tmp_Control_Array(193));
    Control_Array194 <= std_logic_vector(tmp_Control_Array(194));
    Control_Array195 <= std_logic_vector(tmp_Control_Array(195));
    Control_Array196 <= std_logic_vector(tmp_Control_Array(196));
    Control_Array197 <= std_logic_vector(tmp_Control_Array(197));
    Control_Array198 <= std_logic_vector(tmp_Control_Array(198));
    Control_Array199 <= std_logic_vector(tmp_Control_Array(199));
    Control_Array200 <= std_logic_vector(tmp_Control_Array(200));
    Control_Array201 <= std_logic_vector(tmp_Control_Array(201));
    Control_Array202 <= std_logic_vector(tmp_Control_Array(202));
    Control_Array203 <= std_logic_vector(tmp_Control_Array(203));
    Control_Array204 <= std_logic_vector(tmp_Control_Array(204));
    Control_Array205 <= std_logic_vector(tmp_Control_Array(205));
    Control_Array206 <= std_logic_vector(tmp_Control_Array(206));
    Control_Array207 <= std_logic_vector(tmp_Control_Array(207));
    Control_Array208 <= std_logic_vector(tmp_Control_Array(208));
    Control_Array209 <= std_logic_vector(tmp_Control_Array(209));
    Control_Array210 <= std_logic_vector(tmp_Control_Array(210));
    Control_Array211 <= std_logic_vector(tmp_Control_Array(211));
    Control_Array212 <= std_logic_vector(tmp_Control_Array(212));
    Control_Array213 <= std_logic_vector(tmp_Control_Array(213));
    Control_Array214 <= std_logic_vector(tmp_Control_Array(214));
    Control_Array215 <= std_logic_vector(tmp_Control_Array(215));
    Control_Array216 <= std_logic_vector(tmp_Control_Array(216));
    Control_Array217 <= std_logic_vector(tmp_Control_Array(217));
    Control_Array218 <= std_logic_vector(tmp_Control_Array(218));
    Control_Array219 <= std_logic_vector(tmp_Control_Array(219));
    Control_Array220 <= std_logic_vector(tmp_Control_Array(220));
    Control_Array221 <= std_logic_vector(tmp_Control_Array(221));
    Control_Array222 <= std_logic_vector(tmp_Control_Array(222));
    Control_Array223 <= std_logic_vector(tmp_Control_Array(223));
    Control_Array224 <= std_logic_vector(tmp_Control_Array(224));
    Control_Array225 <= std_logic_vector(tmp_Control_Array(225));
    Control_Array226 <= std_logic_vector(tmp_Control_Array(226));
    Control_Array227 <= std_logic_vector(tmp_Control_Array(227));
    Control_Array228 <= std_logic_vector(tmp_Control_Array(228));
    Control_Array229 <= std_logic_vector(tmp_Control_Array(229));
    Control_Array230 <= std_logic_vector(tmp_Control_Array(230));
    Control_Array231 <= std_logic_vector(tmp_Control_Array(231));
    Control_Array232 <= std_logic_vector(tmp_Control_Array(232));
    Control_Array233 <= std_logic_vector(tmp_Control_Array(233));
    Control_Array234 <= std_logic_vector(tmp_Control_Array(234));
    Control_Array235 <= std_logic_vector(tmp_Control_Array(235));
    Control_Array236 <= std_logic_vector(tmp_Control_Array(236));
    Control_Array237 <= std_logic_vector(tmp_Control_Array(237));
    Control_Array238 <= std_logic_vector(tmp_Control_Array(238));
    Control_Array239 <= std_logic_vector(tmp_Control_Array(239));
    Control_Array240 <= std_logic_vector(tmp_Control_Array(240));
    Control_Array241 <= std_logic_vector(tmp_Control_Array(241));
    Control_Array242 <= std_logic_vector(tmp_Control_Array(242));
    Control_Array243 <= std_logic_vector(tmp_Control_Array(243));
    Control_Array244 <= std_logic_vector(tmp_Control_Array(244));
    Control_Array245 <= std_logic_vector(tmp_Control_Array(245));
    Control_Array246 <= std_logic_vector(tmp_Control_Array(246));
    Control_Array247 <= std_logic_vector(tmp_Control_Array(247));
    Control_Array248 <= std_logic_vector(tmp_Control_Array(248));
    Control_Array249 <= std_logic_vector(tmp_Control_Array(249));
    Control_Array250 <= std_logic_vector(tmp_Control_Array(250));
    Control_Array251 <= std_logic_vector(tmp_Control_Array(251));
    Control_Array252 <= std_logic_vector(tmp_Control_Array(252));
    Control_Array253 <= std_logic_vector(tmp_Control_Array(253));
    Control_Array254 <= std_logic_vector(tmp_Control_Array(254));
    Control_Array255 <= std_logic_vector(tmp_Control_Array(255));
    Control_Array256 <= std_logic_vector(tmp_Control_Array(256));
    Control_Array257 <= std_logic_vector(tmp_Control_Array(257));
    Control_Array258 <= std_logic_vector(tmp_Control_Array(258));
    Control_Array259 <= std_logic_vector(tmp_Control_Array(259));
    Control_Array260 <= std_logic_vector(tmp_Control_Array(260));
    Control_Array261 <= std_logic_vector(tmp_Control_Array(261));
    Control_Array262 <= std_logic_vector(tmp_Control_Array(262));
    Control_Array263 <= std_logic_vector(tmp_Control_Array(263));
    Control_Array264 <= std_logic_vector(tmp_Control_Array(264));
    Control_Array265 <= std_logic_vector(tmp_Control_Array(265));
    Control_Array266 <= std_logic_vector(tmp_Control_Array(266));
    Control_Array267 <= std_logic_vector(tmp_Control_Array(267));
    Control_Array268 <= std_logic_vector(tmp_Control_Array(268));
    Control_Array269 <= std_logic_vector(tmp_Control_Array(269));
    Control_Array270 <= std_logic_vector(tmp_Control_Array(270));
    Control_Array271 <= std_logic_vector(tmp_Control_Array(271));
    Control_Array272 <= std_logic_vector(tmp_Control_Array(272));
    Control_Array273 <= std_logic_vector(tmp_Control_Array(273));
    Control_Array274 <= std_logic_vector(tmp_Control_Array(274));
    Control_Array275 <= std_logic_vector(tmp_Control_Array(275));
    Control_Array276 <= std_logic_vector(tmp_Control_Array(276));
    Control_Array277 <= std_logic_vector(tmp_Control_Array(277));
    Control_Array278 <= std_logic_vector(tmp_Control_Array(278));
    Control_Array279 <= std_logic_vector(tmp_Control_Array(279));
    Control_Array280 <= std_logic_vector(tmp_Control_Array(280));
    Control_Array281 <= std_logic_vector(tmp_Control_Array(281));
    Control_Array282 <= std_logic_vector(tmp_Control_Array(282));
    Control_Array283 <= std_logic_vector(tmp_Control_Array(283));
    Control_Array284 <= std_logic_vector(tmp_Control_Array(284));
    Control_Array285 <= std_logic_vector(tmp_Control_Array(285));
    Control_Array286 <= std_logic_vector(tmp_Control_Array(286));
    Control_Array287 <= std_logic_vector(tmp_Control_Array(287));
    Control_Array288 <= std_logic_vector(tmp_Control_Array(288));
    Control_Array289 <= std_logic_vector(tmp_Control_Array(289));
    Control_Array290 <= std_logic_vector(tmp_Control_Array(290));
    Control_Array291 <= std_logic_vector(tmp_Control_Array(291));
    Control_Array292 <= std_logic_vector(tmp_Control_Array(292));
    Control_Array293 <= std_logic_vector(tmp_Control_Array(293));
    Control_Array294 <= std_logic_vector(tmp_Control_Array(294));
    Control_Array295 <= std_logic_vector(tmp_Control_Array(295));
    Control_Array296 <= std_logic_vector(tmp_Control_Array(296));
    Control_Array297 <= std_logic_vector(tmp_Control_Array(297));
    Control_Array298 <= std_logic_vector(tmp_Control_Array(298));
    Control_Array299 <= std_logic_vector(tmp_Control_Array(299));
    Control_Array300 <= std_logic_vector(tmp_Control_Array(300));
    Control_Array301 <= std_logic_vector(tmp_Control_Array(301));
    Control_Array302 <= std_logic_vector(tmp_Control_Array(302));
    Control_Array303 <= std_logic_vector(tmp_Control_Array(303));
    Control_Array304 <= std_logic_vector(tmp_Control_Array(304));
    Control_Array305 <= std_logic_vector(tmp_Control_Array(305));
    Control_Array306 <= std_logic_vector(tmp_Control_Array(306));
    Control_Array307 <= std_logic_vector(tmp_Control_Array(307));
    Control_Array308 <= std_logic_vector(tmp_Control_Array(308));
    Control_Array309 <= std_logic_vector(tmp_Control_Array(309));
    Control_Array310 <= std_logic_vector(tmp_Control_Array(310));
    Control_Array311 <= std_logic_vector(tmp_Control_Array(311));
    Control_Array312 <= std_logic_vector(tmp_Control_Array(312));
    Control_Array313 <= std_logic_vector(tmp_Control_Array(313));
    Control_Array314 <= std_logic_vector(tmp_Control_Array(314));
    Control_Array315 <= std_logic_vector(tmp_Control_Array(315));
    Control_Array316 <= std_logic_vector(tmp_Control_Array(316));
    Control_Array317 <= std_logic_vector(tmp_Control_Array(317));
    Control_Array318 <= std_logic_vector(tmp_Control_Array(318));
    Control_Array319 <= std_logic_vector(tmp_Control_Array(319));
    Control_Array320 <= std_logic_vector(tmp_Control_Array(320));
    Control_Array321 <= std_logic_vector(tmp_Control_Array(321));
    Control_Array322 <= std_logic_vector(tmp_Control_Array(322));
    Control_Array323 <= std_logic_vector(tmp_Control_Array(323));
    Control_Array324 <= std_logic_vector(tmp_Control_Array(324));
    Control_Array325 <= std_logic_vector(tmp_Control_Array(325));
    Control_Array326 <= std_logic_vector(tmp_Control_Array(326));
    Control_Array327 <= std_logic_vector(tmp_Control_Array(327));
    Control_Array328 <= std_logic_vector(tmp_Control_Array(328));
    Control_Array329 <= std_logic_vector(tmp_Control_Array(329));
    Control_Array330 <= std_logic_vector(tmp_Control_Array(330));
    Control_Array331 <= std_logic_vector(tmp_Control_Array(331));
    Control_Array332 <= std_logic_vector(tmp_Control_Array(332));
    Control_Array333 <= std_logic_vector(tmp_Control_Array(333));
    Control_Array334 <= std_logic_vector(tmp_Control_Array(334));
    Control_Array335 <= std_logic_vector(tmp_Control_Array(335));
    Control_Array336 <= std_logic_vector(tmp_Control_Array(336));
    Control_Array337 <= std_logic_vector(tmp_Control_Array(337));
    Control_Array338 <= std_logic_vector(tmp_Control_Array(338));
    Control_Array339 <= std_logic_vector(tmp_Control_Array(339));
    Control_Array340 <= std_logic_vector(tmp_Control_Array(340));
    Control_Array341 <= std_logic_vector(tmp_Control_Array(341));
    Control_Array342 <= std_logic_vector(tmp_Control_Array(342));
    Control_Array343 <= std_logic_vector(tmp_Control_Array(343));
    Control_Array344 <= std_logic_vector(tmp_Control_Array(344));
    Control_Array345 <= std_logic_vector(tmp_Control_Array(345));
    Control_Array346 <= std_logic_vector(tmp_Control_Array(346));
    Control_Array347 <= std_logic_vector(tmp_Control_Array(347));
    Control_Array348 <= std_logic_vector(tmp_Control_Array(348));
    Control_Array349 <= std_logic_vector(tmp_Control_Array(349));
    Control_Array350 <= std_logic_vector(tmp_Control_Array(350));
    Control_Array351 <= std_logic_vector(tmp_Control_Array(351));
    Control_Array352 <= std_logic_vector(tmp_Control_Array(352));
    Control_Array353 <= std_logic_vector(tmp_Control_Array(353));
    Control_Array354 <= std_logic_vector(tmp_Control_Array(354));
    Control_Array355 <= std_logic_vector(tmp_Control_Array(355));
    Control_Array356 <= std_logic_vector(tmp_Control_Array(356));
    Control_Array357 <= std_logic_vector(tmp_Control_Array(357));
    Control_Array358 <= std_logic_vector(tmp_Control_Array(358));
    Control_Array359 <= std_logic_vector(tmp_Control_Array(359));
    Control_Array360 <= std_logic_vector(tmp_Control_Array(360));
    Control_Array361 <= std_logic_vector(tmp_Control_Array(361));
    Control_Array362 <= std_logic_vector(tmp_Control_Array(362));
    Control_Array363 <= std_logic_vector(tmp_Control_Array(363));
    Control_Array364 <= std_logic_vector(tmp_Control_Array(364));
    Control_Array365 <= std_logic_vector(tmp_Control_Array(365));
    Control_Array366 <= std_logic_vector(tmp_Control_Array(366));
    Control_Array367 <= std_logic_vector(tmp_Control_Array(367));
    Control_Array368 <= std_logic_vector(tmp_Control_Array(368));
    Control_Array369 <= std_logic_vector(tmp_Control_Array(369));
    Control_Array370 <= std_logic_vector(tmp_Control_Array(370));
    Control_Array371 <= std_logic_vector(tmp_Control_Array(371));
    Control_Array372 <= std_logic_vector(tmp_Control_Array(372));
    Control_Array373 <= std_logic_vector(tmp_Control_Array(373));
    Control_Array374 <= std_logic_vector(tmp_Control_Array(374));
    Control_Array375 <= std_logic_vector(tmp_Control_Array(375));
    Control_Array376 <= std_logic_vector(tmp_Control_Array(376));
    Control_Array377 <= std_logic_vector(tmp_Control_Array(377));
    Control_Array378 <= std_logic_vector(tmp_Control_Array(378));
    Control_Array379 <= std_logic_vector(tmp_Control_Array(379));
    Control_Array380 <= std_logic_vector(tmp_Control_Array(380));
    Control_Array381 <= std_logic_vector(tmp_Control_Array(381));
    Control_Array382 <= std_logic_vector(tmp_Control_Array(382));
    Control_Array383 <= std_logic_vector(tmp_Control_Array(383));
    Control_Array384 <= std_logic_vector(tmp_Control_Array(384));
    Control_Array385 <= std_logic_vector(tmp_Control_Array(385));
    Control_Array386 <= std_logic_vector(tmp_Control_Array(386));
    Control_Array387 <= std_logic_vector(tmp_Control_Array(387));
    Control_Array388 <= std_logic_vector(tmp_Control_Array(388));
    Control_Array389 <= std_logic_vector(tmp_Control_Array(389));
    Control_Array390 <= std_logic_vector(tmp_Control_Array(390));
    Control_Array391 <= std_logic_vector(tmp_Control_Array(391));
    Control_Array392 <= std_logic_vector(tmp_Control_Array(392));
    Control_Array393 <= std_logic_vector(tmp_Control_Array(393));
    Control_Array394 <= std_logic_vector(tmp_Control_Array(394));
    Control_Array395 <= std_logic_vector(tmp_Control_Array(395));
    Control_Array396 <= std_logic_vector(tmp_Control_Array(396));
    Control_Array397 <= std_logic_vector(tmp_Control_Array(397));
    Control_Array398 <= std_logic_vector(tmp_Control_Array(398));
    Control_Array399 <= std_logic_vector(tmp_Control_Array(399));
    Control_Array400 <= std_logic_vector(tmp_Control_Array(400));
    Control_Array401 <= std_logic_vector(tmp_Control_Array(401));
    Control_Array402 <= std_logic_vector(tmp_Control_Array(402));
    Control_Array403 <= std_logic_vector(tmp_Control_Array(403));
    Control_Array404 <= std_logic_vector(tmp_Control_Array(404));
    Control_Array405 <= std_logic_vector(tmp_Control_Array(405));
    Control_Array406 <= std_logic_vector(tmp_Control_Array(406));
    Control_Array407 <= std_logic_vector(tmp_Control_Array(407));
    Control_Array408 <= std_logic_vector(tmp_Control_Array(408));
    Control_Array409 <= std_logic_vector(tmp_Control_Array(409));
    Control_Array410 <= std_logic_vector(tmp_Control_Array(410));
    Control_Array411 <= std_logic_vector(tmp_Control_Array(411));
    Control_Array412 <= std_logic_vector(tmp_Control_Array(412));
    Control_Array413 <= std_logic_vector(tmp_Control_Array(413));
    Control_Array414 <= std_logic_vector(tmp_Control_Array(414));
    Control_Array415 <= std_logic_vector(tmp_Control_Array(415));
    Control_Array416 <= std_logic_vector(tmp_Control_Array(416));
    Control_Array417 <= std_logic_vector(tmp_Control_Array(417));
    Control_Array418 <= std_logic_vector(tmp_Control_Array(418));
    Control_Array419 <= std_logic_vector(tmp_Control_Array(419));
    Control_Array420 <= std_logic_vector(tmp_Control_Array(420));
    Control_Array421 <= std_logic_vector(tmp_Control_Array(421));
    Control_Array422 <= std_logic_vector(tmp_Control_Array(422));
    Control_Array423 <= std_logic_vector(tmp_Control_Array(423));
    Control_Array424 <= std_logic_vector(tmp_Control_Array(424));
    Control_Array425 <= std_logic_vector(tmp_Control_Array(425));
    Control_Array426 <= std_logic_vector(tmp_Control_Array(426));
    Control_Array427 <= std_logic_vector(tmp_Control_Array(427));
    Control_Array428 <= std_logic_vector(tmp_Control_Array(428));
    Control_Array429 <= std_logic_vector(tmp_Control_Array(429));
    Control_Array430 <= std_logic_vector(tmp_Control_Array(430));
    Control_Array431 <= std_logic_vector(tmp_Control_Array(431));
    Control_Array432 <= std_logic_vector(tmp_Control_Array(432));
    Control_Array433 <= std_logic_vector(tmp_Control_Array(433));
    Control_Array434 <= std_logic_vector(tmp_Control_Array(434));
    Control_Array435 <= std_logic_vector(tmp_Control_Array(435));
    Control_Array436 <= std_logic_vector(tmp_Control_Array(436));
    Control_Array437 <= std_logic_vector(tmp_Control_Array(437));
    Control_Array438 <= std_logic_vector(tmp_Control_Array(438));
    Control_Array439 <= std_logic_vector(tmp_Control_Array(439));
    Control_Array440 <= std_logic_vector(tmp_Control_Array(440));
    Control_Array441 <= std_logic_vector(tmp_Control_Array(441));
    Control_Array442 <= std_logic_vector(tmp_Control_Array(442));
    Control_Array443 <= std_logic_vector(tmp_Control_Array(443));
    Control_Array444 <= std_logic_vector(tmp_Control_Array(444));
    Control_Array445 <= std_logic_vector(tmp_Control_Array(445));
    Control_Array446 <= std_logic_vector(tmp_Control_Array(446));
    Control_Array447 <= std_logic_vector(tmp_Control_Array(447));
    Control_Array448 <= std_logic_vector(tmp_Control_Array(448));
    Control_Array449 <= std_logic_vector(tmp_Control_Array(449));
    Control_Array450 <= std_logic_vector(tmp_Control_Array(450));
    Control_Array451 <= std_logic_vector(tmp_Control_Array(451));
    Control_Array452 <= std_logic_vector(tmp_Control_Array(452));
    Control_Array453 <= std_logic_vector(tmp_Control_Array(453));
    Control_Array454 <= std_logic_vector(tmp_Control_Array(454));
    Control_Array455 <= std_logic_vector(tmp_Control_Array(455));
    Control_Array456 <= std_logic_vector(tmp_Control_Array(456));
    Control_Array457 <= std_logic_vector(tmp_Control_Array(457));
    Control_Array458 <= std_logic_vector(tmp_Control_Array(458));
    Control_Array459 <= std_logic_vector(tmp_Control_Array(459));
    Control_Array460 <= std_logic_vector(tmp_Control_Array(460));
    Control_Array461 <= std_logic_vector(tmp_Control_Array(461));
    Control_Array462 <= std_logic_vector(tmp_Control_Array(462));
    Control_Array463 <= std_logic_vector(tmp_Control_Array(463));
    Control_Array464 <= std_logic_vector(tmp_Control_Array(464));
    Control_Array465 <= std_logic_vector(tmp_Control_Array(465));
    Control_Array466 <= std_logic_vector(tmp_Control_Array(466));
    Control_Array467 <= std_logic_vector(tmp_Control_Array(467));
    Control_Array468 <= std_logic_vector(tmp_Control_Array(468));
    Control_Array469 <= std_logic_vector(tmp_Control_Array(469));
    Control_Array470 <= std_logic_vector(tmp_Control_Array(470));
    Control_Array471 <= std_logic_vector(tmp_Control_Array(471));
    Control_Array472 <= std_logic_vector(tmp_Control_Array(472));
    Control_Array473 <= std_logic_vector(tmp_Control_Array(473));
    Control_Array474 <= std_logic_vector(tmp_Control_Array(474));
    Control_Array475 <= std_logic_vector(tmp_Control_Array(475));
    Control_Array476 <= std_logic_vector(tmp_Control_Array(476));
    Control_Array477 <= std_logic_vector(tmp_Control_Array(477));
    Control_Array478 <= std_logic_vector(tmp_Control_Array(478));
    Control_Array479 <= std_logic_vector(tmp_Control_Array(479));
    Control_Array480 <= std_logic_vector(tmp_Control_Array(480));
    Control_Array481 <= std_logic_vector(tmp_Control_Array(481));
    Control_Array482 <= std_logic_vector(tmp_Control_Array(482));
    Control_Array483 <= std_logic_vector(tmp_Control_Array(483));
    Control_Array484 <= std_logic_vector(tmp_Control_Array(484));
    Control_Array485 <= std_logic_vector(tmp_Control_Array(485));
    Control_Array486 <= std_logic_vector(tmp_Control_Array(486));
    Control_Array487 <= std_logic_vector(tmp_Control_Array(487));
    Control_Array488 <= std_logic_vector(tmp_Control_Array(488));
    Control_Array489 <= std_logic_vector(tmp_Control_Array(489));
    Control_Array490 <= std_logic_vector(tmp_Control_Array(490));
    Control_Array491 <= std_logic_vector(tmp_Control_Array(491));
    Control_Array492 <= std_logic_vector(tmp_Control_Array(492));
    Control_Array493 <= std_logic_vector(tmp_Control_Array(493));
    Control_Array494 <= std_logic_vector(tmp_Control_Array(494));
    Control_Array495 <= std_logic_vector(tmp_Control_Array(495));
    Control_Array496 <= std_logic_vector(tmp_Control_Array(496));
    Control_Array497 <= std_logic_vector(tmp_Control_Array(497));
    Control_Array498 <= std_logic_vector(tmp_Control_Array(498));
    Control_Array499 <= std_logic_vector(tmp_Control_Array(499));
    Control_Array500 <= std_logic_vector(tmp_Control_Array(500));
    Control_Array501 <= std_logic_vector(tmp_Control_Array(501));
    Control_Array502 <= std_logic_vector(tmp_Control_Array(502));
    Control_Array503 <= std_logic_vector(tmp_Control_Array(503));
    Control_Array504 <= std_logic_vector(tmp_Control_Array(504));
    Control_Array505 <= std_logic_vector(tmp_Control_Array(505));
    Control_Array506 <= std_logic_vector(tmp_Control_Array(506));
    Control_Array507 <= std_logic_vector(tmp_Control_Array(507));
    Control_Array508 <= std_logic_vector(tmp_Control_Array(508));
    Control_Array509 <= std_logic_vector(tmp_Control_Array(509));
    Control_Array510 <= std_logic_vector(tmp_Control_Array(510));
    Control_Array511 <= std_logic_vector(tmp_Control_Array(511));
    Control_Array512 <= std_logic_vector(tmp_Control_Array(512));
    Control_Array513 <= std_logic_vector(tmp_Control_Array(513));
    Control_Array514 <= std_logic_vector(tmp_Control_Array(514));
    Control_Array515 <= std_logic_vector(tmp_Control_Array(515));
    Control_Array516 <= std_logic_vector(tmp_Control_Array(516));
    Control_Array517 <= std_logic_vector(tmp_Control_Array(517));
    Control_Array518 <= std_logic_vector(tmp_Control_Array(518));
    Control_Array519 <= std_logic_vector(tmp_Control_Array(519));
    Control_Array520 <= std_logic_vector(tmp_Control_Array(520));
    Control_Array521 <= std_logic_vector(tmp_Control_Array(521));
    Control_Array522 <= std_logic_vector(tmp_Control_Array(522));
    Control_Array523 <= std_logic_vector(tmp_Control_Array(523));
    Control_Array524 <= std_logic_vector(tmp_Control_Array(524));
    Control_Array525 <= std_logic_vector(tmp_Control_Array(525));
    Control_Array526 <= std_logic_vector(tmp_Control_Array(526));
    Control_Array527 <= std_logic_vector(tmp_Control_Array(527));
    Control_Array528 <= std_logic_vector(tmp_Control_Array(528));
    Control_Array529 <= std_logic_vector(tmp_Control_Array(529));
    Control_Array530 <= std_logic_vector(tmp_Control_Array(530));
    Control_Array531 <= std_logic_vector(tmp_Control_Array(531));
    Control_Array532 <= std_logic_vector(tmp_Control_Array(532));
    Control_Array533 <= std_logic_vector(tmp_Control_Array(533));
    Control_Array534 <= std_logic_vector(tmp_Control_Array(534));
    Control_Array535 <= std_logic_vector(tmp_Control_Array(535));
    Control_Array536 <= std_logic_vector(tmp_Control_Array(536));
    Control_Array537 <= std_logic_vector(tmp_Control_Array(537));
    Control_Array538 <= std_logic_vector(tmp_Control_Array(538));
    Control_Array539 <= std_logic_vector(tmp_Control_Array(539));
    Control_Array540 <= std_logic_vector(tmp_Control_Array(540));
    Control_Array541 <= std_logic_vector(tmp_Control_Array(541));
    Control_Array542 <= std_logic_vector(tmp_Control_Array(542));
    Control_Array543 <= std_logic_vector(tmp_Control_Array(543));
    Control_Array544 <= std_logic_vector(tmp_Control_Array(544));
    Control_Array545 <= std_logic_vector(tmp_Control_Array(545));
    Control_Array546 <= std_logic_vector(tmp_Control_Array(546));
    Control_Array547 <= std_logic_vector(tmp_Control_Array(547));
    Control_Array548 <= std_logic_vector(tmp_Control_Array(548));
    Control_Array549 <= std_logic_vector(tmp_Control_Array(549));
    Control_Array550 <= std_logic_vector(tmp_Control_Array(550));
    Control_Array551 <= std_logic_vector(tmp_Control_Array(551));
    Control_Array552 <= std_logic_vector(tmp_Control_Array(552));
    Control_Array553 <= std_logic_vector(tmp_Control_Array(553));
    Control_Array554 <= std_logic_vector(tmp_Control_Array(554));
    Control_Array555 <= std_logic_vector(tmp_Control_Array(555));
    Control_Array556 <= std_logic_vector(tmp_Control_Array(556));
    Control_Array557 <= std_logic_vector(tmp_Control_Array(557));
    Control_Array558 <= std_logic_vector(tmp_Control_Array(558));
    Control_Array559 <= std_logic_vector(tmp_Control_Array(559));
    Control_Array560 <= std_logic_vector(tmp_Control_Array(560));
    Control_Array561 <= std_logic_vector(tmp_Control_Array(561));
    Control_Array562 <= std_logic_vector(tmp_Control_Array(562));
    Control_Array563 <= std_logic_vector(tmp_Control_Array(563));
    Control_Array564 <= std_logic_vector(tmp_Control_Array(564));
    Control_Array565 <= std_logic_vector(tmp_Control_Array(565));
    Control_Array566 <= std_logic_vector(tmp_Control_Array(566));
    Control_Array567 <= std_logic_vector(tmp_Control_Array(567));
    Control_Array568 <= std_logic_vector(tmp_Control_Array(568));
    Control_Array569 <= std_logic_vector(tmp_Control_Array(569));
    Control_Array570 <= std_logic_vector(tmp_Control_Array(570));
    Control_Array571 <= std_logic_vector(tmp_Control_Array(571));
    Control_Array572 <= std_logic_vector(tmp_Control_Array(572));
    Control_Array573 <= std_logic_vector(tmp_Control_Array(573));
    Control_Array574 <= std_logic_vector(tmp_Control_Array(574));
    Control_Array575 <= std_logic_vector(tmp_Control_Array(575));
    Control_Array576 <= std_logic_vector(tmp_Control_Array(576));
    Control_Array577 <= std_logic_vector(tmp_Control_Array(577));
    Control_Array578 <= std_logic_vector(tmp_Control_Array(578));
    Control_Array579 <= std_logic_vector(tmp_Control_Array(579));
    Control_Array580 <= std_logic_vector(tmp_Control_Array(580));
    Control_Array581 <= std_logic_vector(tmp_Control_Array(581));
    Control_Array582 <= std_logic_vector(tmp_Control_Array(582));
    Control_Array583 <= std_logic_vector(tmp_Control_Array(583));
    Control_Array584 <= std_logic_vector(tmp_Control_Array(584));
    Control_Array585 <= std_logic_vector(tmp_Control_Array(585));
    Control_Array586 <= std_logic_vector(tmp_Control_Array(586));
    Control_Array587 <= std_logic_vector(tmp_Control_Array(587));
    Control_Array588 <= std_logic_vector(tmp_Control_Array(588));
    Control_Array589 <= std_logic_vector(tmp_Control_Array(589));
    Control_Array590 <= std_logic_vector(tmp_Control_Array(590));
    Control_Array591 <= std_logic_vector(tmp_Control_Array(591));
    Control_Array592 <= std_logic_vector(tmp_Control_Array(592));
    Control_Array593 <= std_logic_vector(tmp_Control_Array(593));
    Control_Array594 <= std_logic_vector(tmp_Control_Array(594));
    Control_Array595 <= std_logic_vector(tmp_Control_Array(595));
    Control_Array596 <= std_logic_vector(tmp_Control_Array(596));
    Control_Array597 <= std_logic_vector(tmp_Control_Array(597));
    Control_Array598 <= std_logic_vector(tmp_Control_Array(598));
    Control_Array599 <= std_logic_vector(tmp_Control_Array(599));
    Control_Array600 <= std_logic_vector(tmp_Control_Array(600));
    Control_Array601 <= std_logic_vector(tmp_Control_Array(601));
    Control_Array602 <= std_logic_vector(tmp_Control_Array(602));
    Control_Array603 <= std_logic_vector(tmp_Control_Array(603));
    Control_Array604 <= std_logic_vector(tmp_Control_Array(604));
    Control_Array605 <= std_logic_vector(tmp_Control_Array(605));
    Control_Array606 <= std_logic_vector(tmp_Control_Array(606));
    Control_Array607 <= std_logic_vector(tmp_Control_Array(607));
    Control_Array608 <= std_logic_vector(tmp_Control_Array(608));
    Control_Array609 <= std_logic_vector(tmp_Control_Array(609));
    Control_Array610 <= std_logic_vector(tmp_Control_Array(610));
    Control_Array611 <= std_logic_vector(tmp_Control_Array(611));
    Control_Array612 <= std_logic_vector(tmp_Control_Array(612));
    Control_Array613 <= std_logic_vector(tmp_Control_Array(613));
    Control_Array614 <= std_logic_vector(tmp_Control_Array(614));
    Control_Array615 <= std_logic_vector(tmp_Control_Array(615));
    Control_Array616 <= std_logic_vector(tmp_Control_Array(616));
    Control_Array617 <= std_logic_vector(tmp_Control_Array(617));
    Control_Array618 <= std_logic_vector(tmp_Control_Array(618));
    Control_Array619 <= std_logic_vector(tmp_Control_Array(619));
    Control_Array620 <= std_logic_vector(tmp_Control_Array(620));
    Control_Array621 <= std_logic_vector(tmp_Control_Array(621));
    Control_Array622 <= std_logic_vector(tmp_Control_Array(622));
    Control_Array623 <= std_logic_vector(tmp_Control_Array(623));
    Control_Array624 <= std_logic_vector(tmp_Control_Array(624));
    Control_Array625 <= std_logic_vector(tmp_Control_Array(625));
    Control_Array626 <= std_logic_vector(tmp_Control_Array(626));
    Control_Array627 <= std_logic_vector(tmp_Control_Array(627));
    Control_Array628 <= std_logic_vector(tmp_Control_Array(628));
    Control_Array629 <= std_logic_vector(tmp_Control_Array(629));
    Control_Array630 <= std_logic_vector(tmp_Control_Array(630));
    Control_Array631 <= std_logic_vector(tmp_Control_Array(631));
    Control_Array632 <= std_logic_vector(tmp_Control_Array(632));
    Control_Array633 <= std_logic_vector(tmp_Control_Array(633));
    Control_Array634 <= std_logic_vector(tmp_Control_Array(634));
    Control_Array635 <= std_logic_vector(tmp_Control_Array(635));
    Control_Array636 <= std_logic_vector(tmp_Control_Array(636));
    Control_Array637 <= std_logic_vector(tmp_Control_Array(637));
    Control_Array638 <= std_logic_vector(tmp_Control_Array(638));
    Control_Array639 <= std_logic_vector(tmp_Control_Array(639));
    Control_Array640 <= std_logic_vector(tmp_Control_Array(640));
    Control_Array641 <= std_logic_vector(tmp_Control_Array(641));
    Control_Array642 <= std_logic_vector(tmp_Control_Array(642));
    Control_Array643 <= std_logic_vector(tmp_Control_Array(643));
    Control_Array644 <= std_logic_vector(tmp_Control_Array(644));
    Control_Array645 <= std_logic_vector(tmp_Control_Array(645));
    Control_Array646 <= std_logic_vector(tmp_Control_Array(646));
    Control_Array647 <= std_logic_vector(tmp_Control_Array(647));
    Control_Array648 <= std_logic_vector(tmp_Control_Array(648));
    Control_Array649 <= std_logic_vector(tmp_Control_Array(649));
    Control_Array650 <= std_logic_vector(tmp_Control_Array(650));
    Control_Array651 <= std_logic_vector(tmp_Control_Array(651));
    Control_Array652 <= std_logic_vector(tmp_Control_Array(652));
    Control_Array653 <= std_logic_vector(tmp_Control_Array(653));
    Control_Array654 <= std_logic_vector(tmp_Control_Array(654));
    Control_Array655 <= std_logic_vector(tmp_Control_Array(655));
    Control_Array656 <= std_logic_vector(tmp_Control_Array(656));
    Control_Array657 <= std_logic_vector(tmp_Control_Array(657));
    Control_Array658 <= std_logic_vector(tmp_Control_Array(658));
    Control_Array659 <= std_logic_vector(tmp_Control_Array(659));
    Control_Array660 <= std_logic_vector(tmp_Control_Array(660));
    Control_Array661 <= std_logic_vector(tmp_Control_Array(661));
    Control_Array662 <= std_logic_vector(tmp_Control_Array(662));
    Control_Array663 <= std_logic_vector(tmp_Control_Array(663));
    Control_Array664 <= std_logic_vector(tmp_Control_Array(664));
    Control_Array665 <= std_logic_vector(tmp_Control_Array(665));
    Control_Array666 <= std_logic_vector(tmp_Control_Array(666));
    Control_Array667 <= std_logic_vector(tmp_Control_Array(667));
    Control_Array668 <= std_logic_vector(tmp_Control_Array(668));
    Control_Array669 <= std_logic_vector(tmp_Control_Array(669));
    Control_Array670 <= std_logic_vector(tmp_Control_Array(670));
    Control_Array671 <= std_logic_vector(tmp_Control_Array(671));
    Control_Array672 <= std_logic_vector(tmp_Control_Array(672));
    Control_Array673 <= std_logic_vector(tmp_Control_Array(673));
    Control_Array674 <= std_logic_vector(tmp_Control_Array(674));
    Control_Array675 <= std_logic_vector(tmp_Control_Array(675));
    Control_Array676 <= std_logic_vector(tmp_Control_Array(676));
    Control_Array677 <= std_logic_vector(tmp_Control_Array(677));
    Control_Array678 <= std_logic_vector(tmp_Control_Array(678));
    Control_Array679 <= std_logic_vector(tmp_Control_Array(679));
    Control_Array680 <= std_logic_vector(tmp_Control_Array(680));
    Control_Array681 <= std_logic_vector(tmp_Control_Array(681));
    Control_Array682 <= std_logic_vector(tmp_Control_Array(682));
    Control_Array683 <= std_logic_vector(tmp_Control_Array(683));
    Control_Array684 <= std_logic_vector(tmp_Control_Array(684));
    Control_Array685 <= std_logic_vector(tmp_Control_Array(685));
    Control_Array686 <= std_logic_vector(tmp_Control_Array(686));
    Control_Array687 <= std_logic_vector(tmp_Control_Array(687));
    Control_Array688 <= std_logic_vector(tmp_Control_Array(688));
    Control_Array689 <= std_logic_vector(tmp_Control_Array(689));
    Control_Array690 <= std_logic_vector(tmp_Control_Array(690));
    Control_Array691 <= std_logic_vector(tmp_Control_Array(691));
    Control_Array692 <= std_logic_vector(tmp_Control_Array(692));
    Control_Array693 <= std_logic_vector(tmp_Control_Array(693));
    Control_Array694 <= std_logic_vector(tmp_Control_Array(694));
    Control_Array695 <= std_logic_vector(tmp_Control_Array(695));
    Control_Array696 <= std_logic_vector(tmp_Control_Array(696));
    Control_Array697 <= std_logic_vector(tmp_Control_Array(697));
    Control_Array698 <= std_logic_vector(tmp_Control_Array(698));
    Control_Array699 <= std_logic_vector(tmp_Control_Array(699));
    Control_Array700 <= std_logic_vector(tmp_Control_Array(700));
    Control_Array701 <= std_logic_vector(tmp_Control_Array(701));
    Control_Array702 <= std_logic_vector(tmp_Control_Array(702));
    Control_Array703 <= std_logic_vector(tmp_Control_Array(703));
    Control_Array704 <= std_logic_vector(tmp_Control_Array(704));
    Control_Array705 <= std_logic_vector(tmp_Control_Array(705));
    Control_Array706 <= std_logic_vector(tmp_Control_Array(706));
    Control_Array707 <= std_logic_vector(tmp_Control_Array(707));
    Control_Array708 <= std_logic_vector(tmp_Control_Array(708));
    Control_Array709 <= std_logic_vector(tmp_Control_Array(709));
    Control_Array710 <= std_logic_vector(tmp_Control_Array(710));
    Control_Array711 <= std_logic_vector(tmp_Control_Array(711));
    Control_Array712 <= std_logic_vector(tmp_Control_Array(712));
    Control_Array713 <= std_logic_vector(tmp_Control_Array(713));
    Control_Array714 <= std_logic_vector(tmp_Control_Array(714));
    Control_Array715 <= std_logic_vector(tmp_Control_Array(715));
    Control_Array716 <= std_logic_vector(tmp_Control_Array(716));
    Control_Array717 <= std_logic_vector(tmp_Control_Array(717));
    Control_Array718 <= std_logic_vector(tmp_Control_Array(718));
    Control_Array719 <= std_logic_vector(tmp_Control_Array(719));
    Control_Array720 <= std_logic_vector(tmp_Control_Array(720));
    Control_Array721 <= std_logic_vector(tmp_Control_Array(721));
    Control_Array722 <= std_logic_vector(tmp_Control_Array(722));
    Control_Array723 <= std_logic_vector(tmp_Control_Array(723));
    Control_Array724 <= std_logic_vector(tmp_Control_Array(724));
    Control_Array725 <= std_logic_vector(tmp_Control_Array(725));
    Control_Array726 <= std_logic_vector(tmp_Control_Array(726));
    Control_Array727 <= std_logic_vector(tmp_Control_Array(727));
    Control_Array728 <= std_logic_vector(tmp_Control_Array(728));
    Control_Array729 <= std_logic_vector(tmp_Control_Array(729));
    Control_Array730 <= std_logic_vector(tmp_Control_Array(730));
    Control_Array731 <= std_logic_vector(tmp_Control_Array(731));
    Control_Array732 <= std_logic_vector(tmp_Control_Array(732));
    Control_Array733 <= std_logic_vector(tmp_Control_Array(733));
    Control_Array734 <= std_logic_vector(tmp_Control_Array(734));
    Control_Array735 <= std_logic_vector(tmp_Control_Array(735));
    Control_Array736 <= std_logic_vector(tmp_Control_Array(736));
    Control_Array737 <= std_logic_vector(tmp_Control_Array(737));
    Control_Array738 <= std_logic_vector(tmp_Control_Array(738));
    Control_Array739 <= std_logic_vector(tmp_Control_Array(739));
    Control_Array740 <= std_logic_vector(tmp_Control_Array(740));
    Control_Array741 <= std_logic_vector(tmp_Control_Array(741));
    Control_Array742 <= std_logic_vector(tmp_Control_Array(742));
    Control_Array743 <= std_logic_vector(tmp_Control_Array(743));
    Control_Array744 <= std_logic_vector(tmp_Control_Array(744));
    Control_Array745 <= std_logic_vector(tmp_Control_Array(745));
    Control_Array746 <= std_logic_vector(tmp_Control_Array(746));
    Control_Array747 <= std_logic_vector(tmp_Control_Array(747));
    Control_Array748 <= std_logic_vector(tmp_Control_Array(748));
    Control_Array749 <= std_logic_vector(tmp_Control_Array(749));
    Control_Array750 <= std_logic_vector(tmp_Control_Array(750));
    Control_Array751 <= std_logic_vector(tmp_Control_Array(751));
    Control_Array752 <= std_logic_vector(tmp_Control_Array(752));
    Control_Array753 <= std_logic_vector(tmp_Control_Array(753));
    Control_Array754 <= std_logic_vector(tmp_Control_Array(754));
    Control_Array755 <= std_logic_vector(tmp_Control_Array(755));
    Control_Array756 <= std_logic_vector(tmp_Control_Array(756));
    Control_Array757 <= std_logic_vector(tmp_Control_Array(757));
    Control_Array758 <= std_logic_vector(tmp_Control_Array(758));
    Control_Array759 <= std_logic_vector(tmp_Control_Array(759));
    Control_Array760 <= std_logic_vector(tmp_Control_Array(760));
    Control_Array761 <= std_logic_vector(tmp_Control_Array(761));
    Control_Array762 <= std_logic_vector(tmp_Control_Array(762));
    Control_Array763 <= std_logic_vector(tmp_Control_Array(763));
    Control_Array764 <= std_logic_vector(tmp_Control_Array(764));
    Control_Array765 <= std_logic_vector(tmp_Control_Array(765));
    Control_Array766 <= std_logic_vector(tmp_Control_Array(766));
    Control_Array767 <= std_logic_vector(tmp_Control_Array(767));
    Control_Array768 <= std_logic_vector(tmp_Control_Array(768));
    Control_Array769 <= std_logic_vector(tmp_Control_Array(769));
    Control_Array770 <= std_logic_vector(tmp_Control_Array(770));
    Control_Array771 <= std_logic_vector(tmp_Control_Array(771));
    Control_Array772 <= std_logic_vector(tmp_Control_Array(772));
    Control_Array773 <= std_logic_vector(tmp_Control_Array(773));
    Control_Array774 <= std_logic_vector(tmp_Control_Array(774));
    Control_Array775 <= std_logic_vector(tmp_Control_Array(775));
    Control_Array776 <= std_logic_vector(tmp_Control_Array(776));
    Control_Array777 <= std_logic_vector(tmp_Control_Array(777));
    Control_Array778 <= std_logic_vector(tmp_Control_Array(778));
    Control_Array779 <= std_logic_vector(tmp_Control_Array(779));
    Control_Array780 <= std_logic_vector(tmp_Control_Array(780));
    Control_Array781 <= std_logic_vector(tmp_Control_Array(781));
    Control_Array782 <= std_logic_vector(tmp_Control_Array(782));
    Control_Array783 <= std_logic_vector(tmp_Control_Array(783));
    Control_Array784 <= std_logic_vector(tmp_Control_Array(784));
    Control_Array785 <= std_logic_vector(tmp_Control_Array(785));
    Control_Array786 <= std_logic_vector(tmp_Control_Array(786));
    Control_Array787 <= std_logic_vector(tmp_Control_Array(787));
    Control_Array788 <= std_logic_vector(tmp_Control_Array(788));
    Control_Array789 <= std_logic_vector(tmp_Control_Array(789));
    Control_Array790 <= std_logic_vector(tmp_Control_Array(790));
    Control_Array791 <= std_logic_vector(tmp_Control_Array(791));
    Control_Array792 <= std_logic_vector(tmp_Control_Array(792));
    Control_Array793 <= std_logic_vector(tmp_Control_Array(793));
    Control_Array794 <= std_logic_vector(tmp_Control_Array(794));
    Control_Array795 <= std_logic_vector(tmp_Control_Array(795));
    Control_Array796 <= std_logic_vector(tmp_Control_Array(796));
    Control_Array797 <= std_logic_vector(tmp_Control_Array(797));
    Control_Array798 <= std_logic_vector(tmp_Control_Array(798));
    Control_Array799 <= std_logic_vector(tmp_Control_Array(799));
    Control_Array800 <= std_logic_vector(tmp_Control_Array(800));
    Control_Array801 <= std_logic_vector(tmp_Control_Array(801));
    Control_Array802 <= std_logic_vector(tmp_Control_Array(802));
    Control_Array803 <= std_logic_vector(tmp_Control_Array(803));
    Control_Array804 <= std_logic_vector(tmp_Control_Array(804));
    Control_Array805 <= std_logic_vector(tmp_Control_Array(805));
    Control_Array806 <= std_logic_vector(tmp_Control_Array(806));
    Control_Array807 <= std_logic_vector(tmp_Control_Array(807));
    Control_Array808 <= std_logic_vector(tmp_Control_Array(808));
    Control_Array809 <= std_logic_vector(tmp_Control_Array(809));
    Control_Array810 <= std_logic_vector(tmp_Control_Array(810));
    Control_Array811 <= std_logic_vector(tmp_Control_Array(811));
    Control_Array812 <= std_logic_vector(tmp_Control_Array(812));
    Control_Array813 <= std_logic_vector(tmp_Control_Array(813));
    Control_Array814 <= std_logic_vector(tmp_Control_Array(814));
    Control_Array815 <= std_logic_vector(tmp_Control_Array(815));
    Control_Array816 <= std_logic_vector(tmp_Control_Array(816));
    Control_Array817 <= std_logic_vector(tmp_Control_Array(817));
    Control_Array818 <= std_logic_vector(tmp_Control_Array(818));
    Control_Array819 <= std_logic_vector(tmp_Control_Array(819));
    Control_Array820 <= std_logic_vector(tmp_Control_Array(820));
    Control_Array821 <= std_logic_vector(tmp_Control_Array(821));
    Control_Array822 <= std_logic_vector(tmp_Control_Array(822));
    Control_Array823 <= std_logic_vector(tmp_Control_Array(823));
    Control_Array824 <= std_logic_vector(tmp_Control_Array(824));
    Control_Array825 <= std_logic_vector(tmp_Control_Array(825));
    Control_Array826 <= std_logic_vector(tmp_Control_Array(826));
    Control_Array827 <= std_logic_vector(tmp_Control_Array(827));
    Control_Array828 <= std_logic_vector(tmp_Control_Array(828));
    Control_Array829 <= std_logic_vector(tmp_Control_Array(829));
    Control_Array830 <= std_logic_vector(tmp_Control_Array(830));
    Control_Array831 <= std_logic_vector(tmp_Control_Array(831));
    Control_Array832 <= std_logic_vector(tmp_Control_Array(832));
    Control_Array833 <= std_logic_vector(tmp_Control_Array(833));
    Control_Array834 <= std_logic_vector(tmp_Control_Array(834));
    Control_Array835 <= std_logic_vector(tmp_Control_Array(835));
    Control_Array836 <= std_logic_vector(tmp_Control_Array(836));
    Control_Array837 <= std_logic_vector(tmp_Control_Array(837));
    Control_Array838 <= std_logic_vector(tmp_Control_Array(838));
    Control_Array839 <= std_logic_vector(tmp_Control_Array(839));
    Control_Array840 <= std_logic_vector(tmp_Control_Array(840));
    Control_Array841 <= std_logic_vector(tmp_Control_Array(841));
    Control_Array842 <= std_logic_vector(tmp_Control_Array(842));
    Control_Array843 <= std_logic_vector(tmp_Control_Array(843));
    Control_Array844 <= std_logic_vector(tmp_Control_Array(844));
    Control_Array845 <= std_logic_vector(tmp_Control_Array(845));
    Control_Array846 <= std_logic_vector(tmp_Control_Array(846));
    Control_Array847 <= std_logic_vector(tmp_Control_Array(847));
    Control_Array848 <= std_logic_vector(tmp_Control_Array(848));
    Control_Array849 <= std_logic_vector(tmp_Control_Array(849));
    Control_Array850 <= std_logic_vector(tmp_Control_Array(850));
    Control_Array851 <= std_logic_vector(tmp_Control_Array(851));
    Control_Array852 <= std_logic_vector(tmp_Control_Array(852));
    Control_Array853 <= std_logic_vector(tmp_Control_Array(853));
    Control_Array854 <= std_logic_vector(tmp_Control_Array(854));
    Control_Array855 <= std_logic_vector(tmp_Control_Array(855));
    Control_Array856 <= std_logic_vector(tmp_Control_Array(856));
    Control_Array857 <= std_logic_vector(tmp_Control_Array(857));
    Control_Array858 <= std_logic_vector(tmp_Control_Array(858));
    Control_Array859 <= std_logic_vector(tmp_Control_Array(859));
    Control_Array860 <= std_logic_vector(tmp_Control_Array(860));
    Control_Array861 <= std_logic_vector(tmp_Control_Array(861));
    Control_Array862 <= std_logic_vector(tmp_Control_Array(862));
    Control_Array863 <= std_logic_vector(tmp_Control_Array(863));
    Control_Array864 <= std_logic_vector(tmp_Control_Array(864));
    Control_Array865 <= std_logic_vector(tmp_Control_Array(865));
    Control_Array866 <= std_logic_vector(tmp_Control_Array(866));
    Control_Array867 <= std_logic_vector(tmp_Control_Array(867));
    Control_Array868 <= std_logic_vector(tmp_Control_Array(868));
    Control_Array869 <= std_logic_vector(tmp_Control_Array(869));
    Control_Array870 <= std_logic_vector(tmp_Control_Array(870));
    Control_Array871 <= std_logic_vector(tmp_Control_Array(871));
    Control_Array872 <= std_logic_vector(tmp_Control_Array(872));
    Control_Array873 <= std_logic_vector(tmp_Control_Array(873));
    Control_Array874 <= std_logic_vector(tmp_Control_Array(874));
    Control_Array875 <= std_logic_vector(tmp_Control_Array(875));
    Control_Array876 <= std_logic_vector(tmp_Control_Array(876));
    Control_Array877 <= std_logic_vector(tmp_Control_Array(877));
    Control_Array878 <= std_logic_vector(tmp_Control_Array(878));
    Control_Array879 <= std_logic_vector(tmp_Control_Array(879));
    Control_Array880 <= std_logic_vector(tmp_Control_Array(880));
    Control_Array881 <= std_logic_vector(tmp_Control_Array(881));
    Control_Array882 <= std_logic_vector(tmp_Control_Array(882));
    Control_Array883 <= std_logic_vector(tmp_Control_Array(883));
    Control_Array884 <= std_logic_vector(tmp_Control_Array(884));
    Control_Array885 <= std_logic_vector(tmp_Control_Array(885));
    Control_Array886 <= std_logic_vector(tmp_Control_Array(886));
    Control_Array887 <= std_logic_vector(tmp_Control_Array(887));
    Control_Array888 <= std_logic_vector(tmp_Control_Array(888));
    Control_Array889 <= std_logic_vector(tmp_Control_Array(889));
    Control_Array890 <= std_logic_vector(tmp_Control_Array(890));
    Control_Array891 <= std_logic_vector(tmp_Control_Array(891));
    Control_Array892 <= std_logic_vector(tmp_Control_Array(892));
    Control_Array893 <= std_logic_vector(tmp_Control_Array(893));
    Control_Array894 <= std_logic_vector(tmp_Control_Array(894));
    Control_Array895 <= std_logic_vector(tmp_Control_Array(895));
    Control_Array896 <= std_logic_vector(tmp_Control_Array(896));
    Control_Array897 <= std_logic_vector(tmp_Control_Array(897));
    Control_Array898 <= std_logic_vector(tmp_Control_Array(898));
    Control_Array899 <= std_logic_vector(tmp_Control_Array(899));
    Control_Array900 <= std_logic_vector(tmp_Control_Array(900));
    Control_Array901 <= std_logic_vector(tmp_Control_Array(901));
    Control_Array902 <= std_logic_vector(tmp_Control_Array(902));
    Control_Array903 <= std_logic_vector(tmp_Control_Array(903));
    Control_Array904 <= std_logic_vector(tmp_Control_Array(904));
    Control_Array905 <= std_logic_vector(tmp_Control_Array(905));
    Control_Array906 <= std_logic_vector(tmp_Control_Array(906));
    Control_Array907 <= std_logic_vector(tmp_Control_Array(907));
    Control_Array908 <= std_logic_vector(tmp_Control_Array(908));
    Control_Array909 <= std_logic_vector(tmp_Control_Array(909));
    Control_Array910 <= std_logic_vector(tmp_Control_Array(910));
    Control_Array911 <= std_logic_vector(tmp_Control_Array(911));
    Control_Array912 <= std_logic_vector(tmp_Control_Array(912));
    Control_Array913 <= std_logic_vector(tmp_Control_Array(913));
    Control_Array914 <= std_logic_vector(tmp_Control_Array(914));
    Control_Array915 <= std_logic_vector(tmp_Control_Array(915));
    Control_Array916 <= std_logic_vector(tmp_Control_Array(916));
    Control_Array917 <= std_logic_vector(tmp_Control_Array(917));
    Control_Array918 <= std_logic_vector(tmp_Control_Array(918));
    Control_Array919 <= std_logic_vector(tmp_Control_Array(919));
    Control_Array920 <= std_logic_vector(tmp_Control_Array(920));
    Control_Array921 <= std_logic_vector(tmp_Control_Array(921));
    Control_Array922 <= std_logic_vector(tmp_Control_Array(922));
    Control_Array923 <= std_logic_vector(tmp_Control_Array(923));
    Control_Array924 <= std_logic_vector(tmp_Control_Array(924));
    Control_Array925 <= std_logic_vector(tmp_Control_Array(925));
    Control_Array926 <= std_logic_vector(tmp_Control_Array(926));
    Control_Array927 <= std_logic_vector(tmp_Control_Array(927));
    Control_Array928 <= std_logic_vector(tmp_Control_Array(928));
    Control_Array929 <= std_logic_vector(tmp_Control_Array(929));
    Control_Array930 <= std_logic_vector(tmp_Control_Array(930));
    Control_Array931 <= std_logic_vector(tmp_Control_Array(931));
    Control_Array932 <= std_logic_vector(tmp_Control_Array(932));
    Control_Array933 <= std_logic_vector(tmp_Control_Array(933));
    Control_Array934 <= std_logic_vector(tmp_Control_Array(934));
    Control_Array935 <= std_logic_vector(tmp_Control_Array(935));
    Control_Array936 <= std_logic_vector(tmp_Control_Array(936));
    Control_Array937 <= std_logic_vector(tmp_Control_Array(937));
    Control_Array938 <= std_logic_vector(tmp_Control_Array(938));
    Control_Array939 <= std_logic_vector(tmp_Control_Array(939));
    Control_Array940 <= std_logic_vector(tmp_Control_Array(940));
    Control_Array941 <= std_logic_vector(tmp_Control_Array(941));
    Control_Array942 <= std_logic_vector(tmp_Control_Array(942));
    Control_Array943 <= std_logic_vector(tmp_Control_Array(943));
    Control_Array944 <= std_logic_vector(tmp_Control_Array(944));
    Control_Array945 <= std_logic_vector(tmp_Control_Array(945));
    Control_Array946 <= std_logic_vector(tmp_Control_Array(946));
    Control_Array947 <= std_logic_vector(tmp_Control_Array(947));
    Control_Array948 <= std_logic_vector(tmp_Control_Array(948));
    Control_Array949 <= std_logic_vector(tmp_Control_Array(949));
    Control_Array950 <= std_logic_vector(tmp_Control_Array(950));
    Control_Array951 <= std_logic_vector(tmp_Control_Array(951));
    Control_Array952 <= std_logic_vector(tmp_Control_Array(952));
    Control_Array953 <= std_logic_vector(tmp_Control_Array(953));
    Control_Array954 <= std_logic_vector(tmp_Control_Array(954));
    Control_Array955 <= std_logic_vector(tmp_Control_Array(955));
    Control_Array956 <= std_logic_vector(tmp_Control_Array(956));
    Control_Array957 <= std_logic_vector(tmp_Control_Array(957));
    Control_Array958 <= std_logic_vector(tmp_Control_Array(958));
    Control_Array959 <= std_logic_vector(tmp_Control_Array(959));
    Control_Array960 <= std_logic_vector(tmp_Control_Array(960));
    Control_Array961 <= std_logic_vector(tmp_Control_Array(961));
    Control_Array962 <= std_logic_vector(tmp_Control_Array(962));
    Control_Array963 <= std_logic_vector(tmp_Control_Array(963));
    Control_Array964 <= std_logic_vector(tmp_Control_Array(964));
    Control_Array965 <= std_logic_vector(tmp_Control_Array(965));
    Control_Array966 <= std_logic_vector(tmp_Control_Array(966));
    Control_Array967 <= std_logic_vector(tmp_Control_Array(967));
    Control_Array968 <= std_logic_vector(tmp_Control_Array(968));
    Control_Array969 <= std_logic_vector(tmp_Control_Array(969));
    Control_Array970 <= std_logic_vector(tmp_Control_Array(970));
    Control_Array971 <= std_logic_vector(tmp_Control_Array(971));
    Control_Array972 <= std_logic_vector(tmp_Control_Array(972));
    Control_Array973 <= std_logic_vector(tmp_Control_Array(973));
    Control_Array974 <= std_logic_vector(tmp_Control_Array(974));
    Control_Array975 <= std_logic_vector(tmp_Control_Array(975));
    Control_Array976 <= std_logic_vector(tmp_Control_Array(976));
    Control_Array977 <= std_logic_vector(tmp_Control_Array(977));
    Control_Array978 <= std_logic_vector(tmp_Control_Array(978));
    Control_Array979 <= std_logic_vector(tmp_Control_Array(979));
    Control_Array980 <= std_logic_vector(tmp_Control_Array(980));
    Control_Array981 <= std_logic_vector(tmp_Control_Array(981));
    Control_Array982 <= std_logic_vector(tmp_Control_Array(982));
    Control_Array983 <= std_logic_vector(tmp_Control_Array(983));
    Control_Array984 <= std_logic_vector(tmp_Control_Array(984));
    Control_Array985 <= std_logic_vector(tmp_Control_Array(985));
    Control_Array986 <= std_logic_vector(tmp_Control_Array(986));
    Control_Array987 <= std_logic_vector(tmp_Control_Array(987));
    Control_Array988 <= std_logic_vector(tmp_Control_Array(988));
    Control_Array989 <= std_logic_vector(tmp_Control_Array(989));
    Control_Array990 <= std_logic_vector(tmp_Control_Array(990));
    Control_Array991 <= std_logic_vector(tmp_Control_Array(991));
    Control_Array992 <= std_logic_vector(tmp_Control_Array(992));
    Control_Array993 <= std_logic_vector(tmp_Control_Array(993));
    Control_Array994 <= std_logic_vector(tmp_Control_Array(994));
    Control_Array995 <= std_logic_vector(tmp_Control_Array(995));
    Control_Array996 <= std_logic_vector(tmp_Control_Array(996));
    Control_Array997 <= std_logic_vector(tmp_Control_Array(997));
    Control_Array998 <= std_logic_vector(tmp_Control_Array(998));
    Control_Array999 <= std_logic_vector(tmp_Control_Array(999));

    -- Entity sme_intro signals
    sme_intro: entity work.sme_intro
    port map (
        -- Output bus Control
        Control_Valid => Control_Valid,
        Control_Reset => Control_Reset,
        Control_Length => tmp_Control_Length,
        Control_Array => tmp_Control_Array,

        -- Input bus Traversal
        Traversal_Valid => Traversal_Valid,

        ENB => ENB,
        RST => RST,
        FIN => FIN,
        CLK => CLK
    );

-- User defined processes here
-- #### USER-DATA-CODE-START
-- #### USER-DATA-CODE-END

end RTL;