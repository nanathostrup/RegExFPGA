library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- library SYSTEM_TYPES;
use work.SYSTEM_TYPES.ALL;

-- library CUSTOM_TYPES;
use work.CUSTOM_TYPES.ALL;

-- User defined packages here
-- #### USER-DATA-IMPORTS-START
-- #### USER-DATA-IMPORTS-END

entity sme_intro_export is
    port(
        -- Top-level bus Control signals
        Control_Valid: in STD_LOGIC;
        Control_Reset: in STD_LOGIC;
        Control_Length: in STD_LOGIC_VECTOR(31 downto 0);
        Control_Array0: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array1: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array2: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array3: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array4: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array5: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array6: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array7: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array8: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array9: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array10: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array11: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array12: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array13: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array14: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array15: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array16: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array17: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array18: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array19: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array20: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array21: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array22: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array23: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array24: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array25: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array26: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array27: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array28: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array29: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array30: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array31: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array32: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array33: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array34: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array35: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array36: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array37: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array38: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array39: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array40: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array41: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array42: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array43: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array44: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array45: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array46: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array47: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array48: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array49: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array50: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array51: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array52: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array53: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array54: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array55: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array56: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array57: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array58: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array59: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array60: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array61: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array62: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array63: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array64: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array65: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array66: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array67: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array68: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array69: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array70: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array71: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array72: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array73: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array74: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array75: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array76: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array77: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array78: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array79: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array80: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array81: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array82: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array83: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array84: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array85: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array86: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array87: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array88: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array89: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array90: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array91: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array92: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array93: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array94: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array95: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array96: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array97: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array98: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array99: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array100: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array101: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array102: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array103: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array104: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array105: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array106: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array107: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array108: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array109: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array110: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array111: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array112: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array113: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array114: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array115: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array116: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array117: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array118: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array119: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array120: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array121: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array122: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array123: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array124: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array125: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array126: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array127: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array128: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array129: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array130: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array131: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array132: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array133: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array134: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array135: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array136: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array137: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array138: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array139: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array140: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array141: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array142: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array143: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array144: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array145: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array146: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array147: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array148: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array149: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array150: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array151: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array152: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array153: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array154: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array155: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array156: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array157: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array158: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array159: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array160: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array161: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array162: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array163: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array164: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array165: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array166: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array167: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array168: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array169: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array170: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array171: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array172: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array173: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array174: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array175: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array176: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array177: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array178: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array179: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array180: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array181: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array182: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array183: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array184: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array185: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array186: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array187: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array188: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array189: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array190: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array191: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array192: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array193: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array194: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array195: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array196: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array197: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array198: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array199: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array200: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array201: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array202: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array203: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array204: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array205: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array206: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array207: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array208: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array209: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array210: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array211: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array212: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array213: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array214: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array215: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array216: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array217: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array218: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array219: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array220: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array221: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array222: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array223: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array224: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array225: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array226: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array227: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array228: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array229: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array230: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array231: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array232: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array233: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array234: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array235: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array236: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array237: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array238: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array239: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array240: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array241: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array242: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array243: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array244: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array245: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array246: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array247: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array248: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array249: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array250: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array251: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array252: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array253: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array254: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array255: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array256: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array257: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array258: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array259: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array260: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array261: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array262: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array263: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array264: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array265: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array266: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array267: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array268: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array269: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array270: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array271: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array272: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array273: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array274: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array275: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array276: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array277: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array278: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array279: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array280: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array281: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array282: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array283: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array284: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array285: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array286: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array287: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array288: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array289: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array290: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array291: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array292: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array293: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array294: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array295: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array296: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array297: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array298: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array299: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array300: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array301: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array302: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array303: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array304: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array305: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array306: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array307: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array308: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array309: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array310: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array311: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array312: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array313: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array314: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array315: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array316: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array317: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array318: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array319: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array320: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array321: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array322: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array323: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array324: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array325: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array326: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array327: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array328: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array329: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array330: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array331: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array332: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array333: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array334: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array335: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array336: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array337: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array338: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array339: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array340: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array341: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array342: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array343: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array344: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array345: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array346: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array347: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array348: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array349: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array350: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array351: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array352: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array353: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array354: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array355: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array356: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array357: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array358: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array359: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array360: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array361: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array362: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array363: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array364: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array365: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array366: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array367: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array368: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array369: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array370: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array371: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array372: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array373: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array374: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array375: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array376: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array377: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array378: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array379: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array380: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array381: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array382: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array383: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array384: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array385: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array386: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array387: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array388: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array389: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array390: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array391: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array392: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array393: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array394: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array395: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array396: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array397: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array398: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array399: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array400: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array401: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array402: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array403: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array404: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array405: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array406: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array407: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array408: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array409: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array410: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array411: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array412: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array413: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array414: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array415: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array416: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array417: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array418: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array419: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array420: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array421: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array422: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array423: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array424: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array425: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array426: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array427: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array428: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array429: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array430: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array431: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array432: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array433: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array434: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array435: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array436: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array437: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array438: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array439: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array440: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array441: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array442: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array443: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array444: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array445: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array446: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array447: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array448: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array449: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array450: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array451: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array452: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array453: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array454: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array455: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array456: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array457: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array458: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array459: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array460: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array461: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array462: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array463: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array464: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array465: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array466: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array467: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array468: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array469: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array470: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array471: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array472: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array473: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array474: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array475: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array476: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array477: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array478: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array479: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array480: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array481: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array482: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array483: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array484: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array485: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array486: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array487: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array488: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array489: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array490: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array491: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array492: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array493: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array494: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array495: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array496: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array497: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array498: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array499: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array500: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array501: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array502: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array503: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array504: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array505: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array506: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array507: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array508: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array509: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array510: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array511: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array512: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array513: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array514: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array515: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array516: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array517: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array518: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array519: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array520: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array521: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array522: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array523: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array524: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array525: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array526: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array527: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array528: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array529: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array530: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array531: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array532: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array533: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array534: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array535: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array536: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array537: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array538: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array539: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array540: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array541: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array542: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array543: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array544: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array545: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array546: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array547: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array548: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array549: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array550: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array551: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array552: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array553: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array554: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array555: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array556: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array557: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array558: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array559: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array560: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array561: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array562: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array563: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array564: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array565: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array566: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array567: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array568: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array569: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array570: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array571: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array572: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array573: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array574: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array575: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array576: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array577: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array578: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array579: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array580: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array581: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array582: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array583: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array584: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array585: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array586: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array587: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array588: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array589: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array590: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array591: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array592: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array593: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array594: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array595: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array596: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array597: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array598: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array599: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array600: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array601: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array602: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array603: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array604: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array605: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array606: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array607: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array608: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array609: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array610: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array611: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array612: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array613: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array614: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array615: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array616: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array617: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array618: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array619: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array620: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array621: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array622: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array623: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array624: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array625: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array626: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array627: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array628: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array629: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array630: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array631: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array632: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array633: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array634: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array635: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array636: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array637: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array638: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array639: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array640: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array641: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array642: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array643: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array644: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array645: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array646: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array647: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array648: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array649: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array650: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array651: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array652: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array653: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array654: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array655: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array656: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array657: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array658: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array659: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array660: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array661: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array662: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array663: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array664: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array665: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array666: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array667: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array668: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array669: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array670: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array671: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array672: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array673: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array674: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array675: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array676: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array677: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array678: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array679: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array680: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array681: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array682: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array683: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array684: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array685: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array686: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array687: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array688: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array689: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array690: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array691: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array692: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array693: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array694: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array695: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array696: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array697: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array698: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array699: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array700: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array701: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array702: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array703: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array704: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array705: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array706: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array707: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array708: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array709: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array710: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array711: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array712: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array713: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array714: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array715: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array716: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array717: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array718: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array719: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array720: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array721: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array722: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array723: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array724: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array725: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array726: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array727: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array728: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array729: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array730: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array731: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array732: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array733: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array734: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array735: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array736: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array737: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array738: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array739: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array740: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array741: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array742: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array743: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array744: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array745: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array746: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array747: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array748: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array749: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array750: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array751: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array752: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array753: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array754: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array755: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array756: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array757: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array758: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array759: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array760: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array761: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array762: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array763: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array764: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array765: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array766: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array767: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array768: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array769: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array770: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array771: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array772: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array773: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array774: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array775: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array776: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array777: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array778: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array779: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array780: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array781: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array782: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array783: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array784: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array785: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array786: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array787: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array788: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array789: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array790: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array791: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array792: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array793: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array794: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array795: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array796: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array797: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array798: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array799: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array800: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array801: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array802: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array803: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array804: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array805: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array806: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array807: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array808: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array809: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array810: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array811: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array812: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array813: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array814: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array815: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array816: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array817: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array818: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array819: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array820: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array821: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array822: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array823: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array824: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array825: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array826: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array827: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array828: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array829: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array830: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array831: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array832: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array833: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array834: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array835: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array836: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array837: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array838: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array839: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array840: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array841: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array842: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array843: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array844: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array845: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array846: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array847: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array848: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array849: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array850: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array851: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array852: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array853: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array854: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array855: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array856: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array857: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array858: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array859: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array860: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array861: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array862: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array863: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array864: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array865: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array866: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array867: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array868: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array869: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array870: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array871: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array872: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array873: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array874: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array875: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array876: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array877: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array878: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array879: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array880: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array881: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array882: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array883: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array884: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array885: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array886: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array887: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array888: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array889: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array890: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array891: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array892: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array893: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array894: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array895: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array896: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array897: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array898: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array899: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array900: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array901: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array902: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array903: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array904: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array905: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array906: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array907: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array908: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array909: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array910: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array911: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array912: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array913: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array914: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array915: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array916: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array917: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array918: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array919: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array920: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array921: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array922: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array923: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array924: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array925: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array926: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array927: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array928: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array929: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array930: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array931: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array932: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array933: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array934: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array935: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array936: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array937: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array938: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array939: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array940: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array941: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array942: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array943: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array944: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array945: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array946: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array947: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array948: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array949: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array950: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array951: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array952: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array953: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array954: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array955: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array956: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array957: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array958: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array959: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array960: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array961: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array962: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array963: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array964: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array965: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array966: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array967: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array968: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array969: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array970: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array971: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array972: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array973: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array974: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array975: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array976: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array977: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array978: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array979: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array980: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array981: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array982: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array983: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array984: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array985: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array986: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array987: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array988: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array989: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array990: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array991: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array992: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array993: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array994: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array995: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array996: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array997: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array998: in STD_LOGIC_VECTOR(7 downto 0);
        Control_Array999: in STD_LOGIC_VECTOR(7 downto 0);

        -- Top-level bus Traversal signals
        Traversal_Valid: out STD_LOGIC;

        -- User defined signals here
        -- #### USER-DATA-ENTITYSIGNALS-START
        -- #### USER-DATA-ENTITYSIGNALS-END

        -- Enable signal
        ENB : in STD_LOGIC;

        -- Reset signal
        RST : in STD_LOGIC;

        -- Finished signal
        FIN : out Std_logic;

        -- Clock signal
        CLK : in STD_LOGIC
    );
end sme_intro_export;

architecture RTL of sme_intro_export is

    -- User defined signals here
    -- #### USER-DATA-SIGNALS-START
    -- #### USER-DATA-SIGNALS-END

    -- Intermediate conversion signal to convert internal types to external ones
    signal tmp_Control_Array : Control_Array_type;

begin

    -- Carry converted signals from entity to wrapped outputs
    tmp_Control_Array(0) <= unsigned(Control_Array0);
    tmp_Control_Array(1) <= unsigned(Control_Array1);
    tmp_Control_Array(2) <= unsigned(Control_Array2);
    tmp_Control_Array(3) <= unsigned(Control_Array3);
    tmp_Control_Array(4) <= unsigned(Control_Array4);
    tmp_Control_Array(5) <= unsigned(Control_Array5);
    tmp_Control_Array(6) <= unsigned(Control_Array6);
    tmp_Control_Array(7) <= unsigned(Control_Array7);
    tmp_Control_Array(8) <= unsigned(Control_Array8);
    tmp_Control_Array(9) <= unsigned(Control_Array9);
    tmp_Control_Array(10) <= unsigned(Control_Array10);
    tmp_Control_Array(11) <= unsigned(Control_Array11);
    tmp_Control_Array(12) <= unsigned(Control_Array12);
    tmp_Control_Array(13) <= unsigned(Control_Array13);
    tmp_Control_Array(14) <= unsigned(Control_Array14);
    tmp_Control_Array(15) <= unsigned(Control_Array15);
    tmp_Control_Array(16) <= unsigned(Control_Array16);
    tmp_Control_Array(17) <= unsigned(Control_Array17);
    tmp_Control_Array(18) <= unsigned(Control_Array18);
    tmp_Control_Array(19) <= unsigned(Control_Array19);
    tmp_Control_Array(20) <= unsigned(Control_Array20);
    tmp_Control_Array(21) <= unsigned(Control_Array21);
    tmp_Control_Array(22) <= unsigned(Control_Array22);
    tmp_Control_Array(23) <= unsigned(Control_Array23);
    tmp_Control_Array(24) <= unsigned(Control_Array24);
    tmp_Control_Array(25) <= unsigned(Control_Array25);
    tmp_Control_Array(26) <= unsigned(Control_Array26);
    tmp_Control_Array(27) <= unsigned(Control_Array27);
    tmp_Control_Array(28) <= unsigned(Control_Array28);
    tmp_Control_Array(29) <= unsigned(Control_Array29);
    tmp_Control_Array(30) <= unsigned(Control_Array30);
    tmp_Control_Array(31) <= unsigned(Control_Array31);
    tmp_Control_Array(32) <= unsigned(Control_Array32);
    tmp_Control_Array(33) <= unsigned(Control_Array33);
    tmp_Control_Array(34) <= unsigned(Control_Array34);
    tmp_Control_Array(35) <= unsigned(Control_Array35);
    tmp_Control_Array(36) <= unsigned(Control_Array36);
    tmp_Control_Array(37) <= unsigned(Control_Array37);
    tmp_Control_Array(38) <= unsigned(Control_Array38);
    tmp_Control_Array(39) <= unsigned(Control_Array39);
    tmp_Control_Array(40) <= unsigned(Control_Array40);
    tmp_Control_Array(41) <= unsigned(Control_Array41);
    tmp_Control_Array(42) <= unsigned(Control_Array42);
    tmp_Control_Array(43) <= unsigned(Control_Array43);
    tmp_Control_Array(44) <= unsigned(Control_Array44);
    tmp_Control_Array(45) <= unsigned(Control_Array45);
    tmp_Control_Array(46) <= unsigned(Control_Array46);
    tmp_Control_Array(47) <= unsigned(Control_Array47);
    tmp_Control_Array(48) <= unsigned(Control_Array48);
    tmp_Control_Array(49) <= unsigned(Control_Array49);
    tmp_Control_Array(50) <= unsigned(Control_Array50);
    tmp_Control_Array(51) <= unsigned(Control_Array51);
    tmp_Control_Array(52) <= unsigned(Control_Array52);
    tmp_Control_Array(53) <= unsigned(Control_Array53);
    tmp_Control_Array(54) <= unsigned(Control_Array54);
    tmp_Control_Array(55) <= unsigned(Control_Array55);
    tmp_Control_Array(56) <= unsigned(Control_Array56);
    tmp_Control_Array(57) <= unsigned(Control_Array57);
    tmp_Control_Array(58) <= unsigned(Control_Array58);
    tmp_Control_Array(59) <= unsigned(Control_Array59);
    tmp_Control_Array(60) <= unsigned(Control_Array60);
    tmp_Control_Array(61) <= unsigned(Control_Array61);
    tmp_Control_Array(62) <= unsigned(Control_Array62);
    tmp_Control_Array(63) <= unsigned(Control_Array63);
    tmp_Control_Array(64) <= unsigned(Control_Array64);
    tmp_Control_Array(65) <= unsigned(Control_Array65);
    tmp_Control_Array(66) <= unsigned(Control_Array66);
    tmp_Control_Array(67) <= unsigned(Control_Array67);
    tmp_Control_Array(68) <= unsigned(Control_Array68);
    tmp_Control_Array(69) <= unsigned(Control_Array69);
    tmp_Control_Array(70) <= unsigned(Control_Array70);
    tmp_Control_Array(71) <= unsigned(Control_Array71);
    tmp_Control_Array(72) <= unsigned(Control_Array72);
    tmp_Control_Array(73) <= unsigned(Control_Array73);
    tmp_Control_Array(74) <= unsigned(Control_Array74);
    tmp_Control_Array(75) <= unsigned(Control_Array75);
    tmp_Control_Array(76) <= unsigned(Control_Array76);
    tmp_Control_Array(77) <= unsigned(Control_Array77);
    tmp_Control_Array(78) <= unsigned(Control_Array78);
    tmp_Control_Array(79) <= unsigned(Control_Array79);
    tmp_Control_Array(80) <= unsigned(Control_Array80);
    tmp_Control_Array(81) <= unsigned(Control_Array81);
    tmp_Control_Array(82) <= unsigned(Control_Array82);
    tmp_Control_Array(83) <= unsigned(Control_Array83);
    tmp_Control_Array(84) <= unsigned(Control_Array84);
    tmp_Control_Array(85) <= unsigned(Control_Array85);
    tmp_Control_Array(86) <= unsigned(Control_Array86);
    tmp_Control_Array(87) <= unsigned(Control_Array87);
    tmp_Control_Array(88) <= unsigned(Control_Array88);
    tmp_Control_Array(89) <= unsigned(Control_Array89);
    tmp_Control_Array(90) <= unsigned(Control_Array90);
    tmp_Control_Array(91) <= unsigned(Control_Array91);
    tmp_Control_Array(92) <= unsigned(Control_Array92);
    tmp_Control_Array(93) <= unsigned(Control_Array93);
    tmp_Control_Array(94) <= unsigned(Control_Array94);
    tmp_Control_Array(95) <= unsigned(Control_Array95);
    tmp_Control_Array(96) <= unsigned(Control_Array96);
    tmp_Control_Array(97) <= unsigned(Control_Array97);
    tmp_Control_Array(98) <= unsigned(Control_Array98);
    tmp_Control_Array(99) <= unsigned(Control_Array99);
    tmp_Control_Array(100) <= unsigned(Control_Array100);
    tmp_Control_Array(101) <= unsigned(Control_Array101);
    tmp_Control_Array(102) <= unsigned(Control_Array102);
    tmp_Control_Array(103) <= unsigned(Control_Array103);
    tmp_Control_Array(104) <= unsigned(Control_Array104);
    tmp_Control_Array(105) <= unsigned(Control_Array105);
    tmp_Control_Array(106) <= unsigned(Control_Array106);
    tmp_Control_Array(107) <= unsigned(Control_Array107);
    tmp_Control_Array(108) <= unsigned(Control_Array108);
    tmp_Control_Array(109) <= unsigned(Control_Array109);
    tmp_Control_Array(110) <= unsigned(Control_Array110);
    tmp_Control_Array(111) <= unsigned(Control_Array111);
    tmp_Control_Array(112) <= unsigned(Control_Array112);
    tmp_Control_Array(113) <= unsigned(Control_Array113);
    tmp_Control_Array(114) <= unsigned(Control_Array114);
    tmp_Control_Array(115) <= unsigned(Control_Array115);
    tmp_Control_Array(116) <= unsigned(Control_Array116);
    tmp_Control_Array(117) <= unsigned(Control_Array117);
    tmp_Control_Array(118) <= unsigned(Control_Array118);
    tmp_Control_Array(119) <= unsigned(Control_Array119);
    tmp_Control_Array(120) <= unsigned(Control_Array120);
    tmp_Control_Array(121) <= unsigned(Control_Array121);
    tmp_Control_Array(122) <= unsigned(Control_Array122);
    tmp_Control_Array(123) <= unsigned(Control_Array123);
    tmp_Control_Array(124) <= unsigned(Control_Array124);
    tmp_Control_Array(125) <= unsigned(Control_Array125);
    tmp_Control_Array(126) <= unsigned(Control_Array126);
    tmp_Control_Array(127) <= unsigned(Control_Array127);
    tmp_Control_Array(128) <= unsigned(Control_Array128);
    tmp_Control_Array(129) <= unsigned(Control_Array129);
    tmp_Control_Array(130) <= unsigned(Control_Array130);
    tmp_Control_Array(131) <= unsigned(Control_Array131);
    tmp_Control_Array(132) <= unsigned(Control_Array132);
    tmp_Control_Array(133) <= unsigned(Control_Array133);
    tmp_Control_Array(134) <= unsigned(Control_Array134);
    tmp_Control_Array(135) <= unsigned(Control_Array135);
    tmp_Control_Array(136) <= unsigned(Control_Array136);
    tmp_Control_Array(137) <= unsigned(Control_Array137);
    tmp_Control_Array(138) <= unsigned(Control_Array138);
    tmp_Control_Array(139) <= unsigned(Control_Array139);
    tmp_Control_Array(140) <= unsigned(Control_Array140);
    tmp_Control_Array(141) <= unsigned(Control_Array141);
    tmp_Control_Array(142) <= unsigned(Control_Array142);
    tmp_Control_Array(143) <= unsigned(Control_Array143);
    tmp_Control_Array(144) <= unsigned(Control_Array144);
    tmp_Control_Array(145) <= unsigned(Control_Array145);
    tmp_Control_Array(146) <= unsigned(Control_Array146);
    tmp_Control_Array(147) <= unsigned(Control_Array147);
    tmp_Control_Array(148) <= unsigned(Control_Array148);
    tmp_Control_Array(149) <= unsigned(Control_Array149);
    tmp_Control_Array(150) <= unsigned(Control_Array150);
    tmp_Control_Array(151) <= unsigned(Control_Array151);
    tmp_Control_Array(152) <= unsigned(Control_Array152);
    tmp_Control_Array(153) <= unsigned(Control_Array153);
    tmp_Control_Array(154) <= unsigned(Control_Array154);
    tmp_Control_Array(155) <= unsigned(Control_Array155);
    tmp_Control_Array(156) <= unsigned(Control_Array156);
    tmp_Control_Array(157) <= unsigned(Control_Array157);
    tmp_Control_Array(158) <= unsigned(Control_Array158);
    tmp_Control_Array(159) <= unsigned(Control_Array159);
    tmp_Control_Array(160) <= unsigned(Control_Array160);
    tmp_Control_Array(161) <= unsigned(Control_Array161);
    tmp_Control_Array(162) <= unsigned(Control_Array162);
    tmp_Control_Array(163) <= unsigned(Control_Array163);
    tmp_Control_Array(164) <= unsigned(Control_Array164);
    tmp_Control_Array(165) <= unsigned(Control_Array165);
    tmp_Control_Array(166) <= unsigned(Control_Array166);
    tmp_Control_Array(167) <= unsigned(Control_Array167);
    tmp_Control_Array(168) <= unsigned(Control_Array168);
    tmp_Control_Array(169) <= unsigned(Control_Array169);
    tmp_Control_Array(170) <= unsigned(Control_Array170);
    tmp_Control_Array(171) <= unsigned(Control_Array171);
    tmp_Control_Array(172) <= unsigned(Control_Array172);
    tmp_Control_Array(173) <= unsigned(Control_Array173);
    tmp_Control_Array(174) <= unsigned(Control_Array174);
    tmp_Control_Array(175) <= unsigned(Control_Array175);
    tmp_Control_Array(176) <= unsigned(Control_Array176);
    tmp_Control_Array(177) <= unsigned(Control_Array177);
    tmp_Control_Array(178) <= unsigned(Control_Array178);
    tmp_Control_Array(179) <= unsigned(Control_Array179);
    tmp_Control_Array(180) <= unsigned(Control_Array180);
    tmp_Control_Array(181) <= unsigned(Control_Array181);
    tmp_Control_Array(182) <= unsigned(Control_Array182);
    tmp_Control_Array(183) <= unsigned(Control_Array183);
    tmp_Control_Array(184) <= unsigned(Control_Array184);
    tmp_Control_Array(185) <= unsigned(Control_Array185);
    tmp_Control_Array(186) <= unsigned(Control_Array186);
    tmp_Control_Array(187) <= unsigned(Control_Array187);
    tmp_Control_Array(188) <= unsigned(Control_Array188);
    tmp_Control_Array(189) <= unsigned(Control_Array189);
    tmp_Control_Array(190) <= unsigned(Control_Array190);
    tmp_Control_Array(191) <= unsigned(Control_Array191);
    tmp_Control_Array(192) <= unsigned(Control_Array192);
    tmp_Control_Array(193) <= unsigned(Control_Array193);
    tmp_Control_Array(194) <= unsigned(Control_Array194);
    tmp_Control_Array(195) <= unsigned(Control_Array195);
    tmp_Control_Array(196) <= unsigned(Control_Array196);
    tmp_Control_Array(197) <= unsigned(Control_Array197);
    tmp_Control_Array(198) <= unsigned(Control_Array198);
    tmp_Control_Array(199) <= unsigned(Control_Array199);
    tmp_Control_Array(200) <= unsigned(Control_Array200);
    tmp_Control_Array(201) <= unsigned(Control_Array201);
    tmp_Control_Array(202) <= unsigned(Control_Array202);
    tmp_Control_Array(203) <= unsigned(Control_Array203);
    tmp_Control_Array(204) <= unsigned(Control_Array204);
    tmp_Control_Array(205) <= unsigned(Control_Array205);
    tmp_Control_Array(206) <= unsigned(Control_Array206);
    tmp_Control_Array(207) <= unsigned(Control_Array207);
    tmp_Control_Array(208) <= unsigned(Control_Array208);
    tmp_Control_Array(209) <= unsigned(Control_Array209);
    tmp_Control_Array(210) <= unsigned(Control_Array210);
    tmp_Control_Array(211) <= unsigned(Control_Array211);
    tmp_Control_Array(212) <= unsigned(Control_Array212);
    tmp_Control_Array(213) <= unsigned(Control_Array213);
    tmp_Control_Array(214) <= unsigned(Control_Array214);
    tmp_Control_Array(215) <= unsigned(Control_Array215);
    tmp_Control_Array(216) <= unsigned(Control_Array216);
    tmp_Control_Array(217) <= unsigned(Control_Array217);
    tmp_Control_Array(218) <= unsigned(Control_Array218);
    tmp_Control_Array(219) <= unsigned(Control_Array219);
    tmp_Control_Array(220) <= unsigned(Control_Array220);
    tmp_Control_Array(221) <= unsigned(Control_Array221);
    tmp_Control_Array(222) <= unsigned(Control_Array222);
    tmp_Control_Array(223) <= unsigned(Control_Array223);
    tmp_Control_Array(224) <= unsigned(Control_Array224);
    tmp_Control_Array(225) <= unsigned(Control_Array225);
    tmp_Control_Array(226) <= unsigned(Control_Array226);
    tmp_Control_Array(227) <= unsigned(Control_Array227);
    tmp_Control_Array(228) <= unsigned(Control_Array228);
    tmp_Control_Array(229) <= unsigned(Control_Array229);
    tmp_Control_Array(230) <= unsigned(Control_Array230);
    tmp_Control_Array(231) <= unsigned(Control_Array231);
    tmp_Control_Array(232) <= unsigned(Control_Array232);
    tmp_Control_Array(233) <= unsigned(Control_Array233);
    tmp_Control_Array(234) <= unsigned(Control_Array234);
    tmp_Control_Array(235) <= unsigned(Control_Array235);
    tmp_Control_Array(236) <= unsigned(Control_Array236);
    tmp_Control_Array(237) <= unsigned(Control_Array237);
    tmp_Control_Array(238) <= unsigned(Control_Array238);
    tmp_Control_Array(239) <= unsigned(Control_Array239);
    tmp_Control_Array(240) <= unsigned(Control_Array240);
    tmp_Control_Array(241) <= unsigned(Control_Array241);
    tmp_Control_Array(242) <= unsigned(Control_Array242);
    tmp_Control_Array(243) <= unsigned(Control_Array243);
    tmp_Control_Array(244) <= unsigned(Control_Array244);
    tmp_Control_Array(245) <= unsigned(Control_Array245);
    tmp_Control_Array(246) <= unsigned(Control_Array246);
    tmp_Control_Array(247) <= unsigned(Control_Array247);
    tmp_Control_Array(248) <= unsigned(Control_Array248);
    tmp_Control_Array(249) <= unsigned(Control_Array249);
    tmp_Control_Array(250) <= unsigned(Control_Array250);
    tmp_Control_Array(251) <= unsigned(Control_Array251);
    tmp_Control_Array(252) <= unsigned(Control_Array252);
    tmp_Control_Array(253) <= unsigned(Control_Array253);
    tmp_Control_Array(254) <= unsigned(Control_Array254);
    tmp_Control_Array(255) <= unsigned(Control_Array255);
    tmp_Control_Array(256) <= unsigned(Control_Array256);
    tmp_Control_Array(257) <= unsigned(Control_Array257);
    tmp_Control_Array(258) <= unsigned(Control_Array258);
    tmp_Control_Array(259) <= unsigned(Control_Array259);
    tmp_Control_Array(260) <= unsigned(Control_Array260);
    tmp_Control_Array(261) <= unsigned(Control_Array261);
    tmp_Control_Array(262) <= unsigned(Control_Array262);
    tmp_Control_Array(263) <= unsigned(Control_Array263);
    tmp_Control_Array(264) <= unsigned(Control_Array264);
    tmp_Control_Array(265) <= unsigned(Control_Array265);
    tmp_Control_Array(266) <= unsigned(Control_Array266);
    tmp_Control_Array(267) <= unsigned(Control_Array267);
    tmp_Control_Array(268) <= unsigned(Control_Array268);
    tmp_Control_Array(269) <= unsigned(Control_Array269);
    tmp_Control_Array(270) <= unsigned(Control_Array270);
    tmp_Control_Array(271) <= unsigned(Control_Array271);
    tmp_Control_Array(272) <= unsigned(Control_Array272);
    tmp_Control_Array(273) <= unsigned(Control_Array273);
    tmp_Control_Array(274) <= unsigned(Control_Array274);
    tmp_Control_Array(275) <= unsigned(Control_Array275);
    tmp_Control_Array(276) <= unsigned(Control_Array276);
    tmp_Control_Array(277) <= unsigned(Control_Array277);
    tmp_Control_Array(278) <= unsigned(Control_Array278);
    tmp_Control_Array(279) <= unsigned(Control_Array279);
    tmp_Control_Array(280) <= unsigned(Control_Array280);
    tmp_Control_Array(281) <= unsigned(Control_Array281);
    tmp_Control_Array(282) <= unsigned(Control_Array282);
    tmp_Control_Array(283) <= unsigned(Control_Array283);
    tmp_Control_Array(284) <= unsigned(Control_Array284);
    tmp_Control_Array(285) <= unsigned(Control_Array285);
    tmp_Control_Array(286) <= unsigned(Control_Array286);
    tmp_Control_Array(287) <= unsigned(Control_Array287);
    tmp_Control_Array(288) <= unsigned(Control_Array288);
    tmp_Control_Array(289) <= unsigned(Control_Array289);
    tmp_Control_Array(290) <= unsigned(Control_Array290);
    tmp_Control_Array(291) <= unsigned(Control_Array291);
    tmp_Control_Array(292) <= unsigned(Control_Array292);
    tmp_Control_Array(293) <= unsigned(Control_Array293);
    tmp_Control_Array(294) <= unsigned(Control_Array294);
    tmp_Control_Array(295) <= unsigned(Control_Array295);
    tmp_Control_Array(296) <= unsigned(Control_Array296);
    tmp_Control_Array(297) <= unsigned(Control_Array297);
    tmp_Control_Array(298) <= unsigned(Control_Array298);
    tmp_Control_Array(299) <= unsigned(Control_Array299);
    tmp_Control_Array(300) <= unsigned(Control_Array300);
    tmp_Control_Array(301) <= unsigned(Control_Array301);
    tmp_Control_Array(302) <= unsigned(Control_Array302);
    tmp_Control_Array(303) <= unsigned(Control_Array303);
    tmp_Control_Array(304) <= unsigned(Control_Array304);
    tmp_Control_Array(305) <= unsigned(Control_Array305);
    tmp_Control_Array(306) <= unsigned(Control_Array306);
    tmp_Control_Array(307) <= unsigned(Control_Array307);
    tmp_Control_Array(308) <= unsigned(Control_Array308);
    tmp_Control_Array(309) <= unsigned(Control_Array309);
    tmp_Control_Array(310) <= unsigned(Control_Array310);
    tmp_Control_Array(311) <= unsigned(Control_Array311);
    tmp_Control_Array(312) <= unsigned(Control_Array312);
    tmp_Control_Array(313) <= unsigned(Control_Array313);
    tmp_Control_Array(314) <= unsigned(Control_Array314);
    tmp_Control_Array(315) <= unsigned(Control_Array315);
    tmp_Control_Array(316) <= unsigned(Control_Array316);
    tmp_Control_Array(317) <= unsigned(Control_Array317);
    tmp_Control_Array(318) <= unsigned(Control_Array318);
    tmp_Control_Array(319) <= unsigned(Control_Array319);
    tmp_Control_Array(320) <= unsigned(Control_Array320);
    tmp_Control_Array(321) <= unsigned(Control_Array321);
    tmp_Control_Array(322) <= unsigned(Control_Array322);
    tmp_Control_Array(323) <= unsigned(Control_Array323);
    tmp_Control_Array(324) <= unsigned(Control_Array324);
    tmp_Control_Array(325) <= unsigned(Control_Array325);
    tmp_Control_Array(326) <= unsigned(Control_Array326);
    tmp_Control_Array(327) <= unsigned(Control_Array327);
    tmp_Control_Array(328) <= unsigned(Control_Array328);
    tmp_Control_Array(329) <= unsigned(Control_Array329);
    tmp_Control_Array(330) <= unsigned(Control_Array330);
    tmp_Control_Array(331) <= unsigned(Control_Array331);
    tmp_Control_Array(332) <= unsigned(Control_Array332);
    tmp_Control_Array(333) <= unsigned(Control_Array333);
    tmp_Control_Array(334) <= unsigned(Control_Array334);
    tmp_Control_Array(335) <= unsigned(Control_Array335);
    tmp_Control_Array(336) <= unsigned(Control_Array336);
    tmp_Control_Array(337) <= unsigned(Control_Array337);
    tmp_Control_Array(338) <= unsigned(Control_Array338);
    tmp_Control_Array(339) <= unsigned(Control_Array339);
    tmp_Control_Array(340) <= unsigned(Control_Array340);
    tmp_Control_Array(341) <= unsigned(Control_Array341);
    tmp_Control_Array(342) <= unsigned(Control_Array342);
    tmp_Control_Array(343) <= unsigned(Control_Array343);
    tmp_Control_Array(344) <= unsigned(Control_Array344);
    tmp_Control_Array(345) <= unsigned(Control_Array345);
    tmp_Control_Array(346) <= unsigned(Control_Array346);
    tmp_Control_Array(347) <= unsigned(Control_Array347);
    tmp_Control_Array(348) <= unsigned(Control_Array348);
    tmp_Control_Array(349) <= unsigned(Control_Array349);
    tmp_Control_Array(350) <= unsigned(Control_Array350);
    tmp_Control_Array(351) <= unsigned(Control_Array351);
    tmp_Control_Array(352) <= unsigned(Control_Array352);
    tmp_Control_Array(353) <= unsigned(Control_Array353);
    tmp_Control_Array(354) <= unsigned(Control_Array354);
    tmp_Control_Array(355) <= unsigned(Control_Array355);
    tmp_Control_Array(356) <= unsigned(Control_Array356);
    tmp_Control_Array(357) <= unsigned(Control_Array357);
    tmp_Control_Array(358) <= unsigned(Control_Array358);
    tmp_Control_Array(359) <= unsigned(Control_Array359);
    tmp_Control_Array(360) <= unsigned(Control_Array360);
    tmp_Control_Array(361) <= unsigned(Control_Array361);
    tmp_Control_Array(362) <= unsigned(Control_Array362);
    tmp_Control_Array(363) <= unsigned(Control_Array363);
    tmp_Control_Array(364) <= unsigned(Control_Array364);
    tmp_Control_Array(365) <= unsigned(Control_Array365);
    tmp_Control_Array(366) <= unsigned(Control_Array366);
    tmp_Control_Array(367) <= unsigned(Control_Array367);
    tmp_Control_Array(368) <= unsigned(Control_Array368);
    tmp_Control_Array(369) <= unsigned(Control_Array369);
    tmp_Control_Array(370) <= unsigned(Control_Array370);
    tmp_Control_Array(371) <= unsigned(Control_Array371);
    tmp_Control_Array(372) <= unsigned(Control_Array372);
    tmp_Control_Array(373) <= unsigned(Control_Array373);
    tmp_Control_Array(374) <= unsigned(Control_Array374);
    tmp_Control_Array(375) <= unsigned(Control_Array375);
    tmp_Control_Array(376) <= unsigned(Control_Array376);
    tmp_Control_Array(377) <= unsigned(Control_Array377);
    tmp_Control_Array(378) <= unsigned(Control_Array378);
    tmp_Control_Array(379) <= unsigned(Control_Array379);
    tmp_Control_Array(380) <= unsigned(Control_Array380);
    tmp_Control_Array(381) <= unsigned(Control_Array381);
    tmp_Control_Array(382) <= unsigned(Control_Array382);
    tmp_Control_Array(383) <= unsigned(Control_Array383);
    tmp_Control_Array(384) <= unsigned(Control_Array384);
    tmp_Control_Array(385) <= unsigned(Control_Array385);
    tmp_Control_Array(386) <= unsigned(Control_Array386);
    tmp_Control_Array(387) <= unsigned(Control_Array387);
    tmp_Control_Array(388) <= unsigned(Control_Array388);
    tmp_Control_Array(389) <= unsigned(Control_Array389);
    tmp_Control_Array(390) <= unsigned(Control_Array390);
    tmp_Control_Array(391) <= unsigned(Control_Array391);
    tmp_Control_Array(392) <= unsigned(Control_Array392);
    tmp_Control_Array(393) <= unsigned(Control_Array393);
    tmp_Control_Array(394) <= unsigned(Control_Array394);
    tmp_Control_Array(395) <= unsigned(Control_Array395);
    tmp_Control_Array(396) <= unsigned(Control_Array396);
    tmp_Control_Array(397) <= unsigned(Control_Array397);
    tmp_Control_Array(398) <= unsigned(Control_Array398);
    tmp_Control_Array(399) <= unsigned(Control_Array399);
    tmp_Control_Array(400) <= unsigned(Control_Array400);
    tmp_Control_Array(401) <= unsigned(Control_Array401);
    tmp_Control_Array(402) <= unsigned(Control_Array402);
    tmp_Control_Array(403) <= unsigned(Control_Array403);
    tmp_Control_Array(404) <= unsigned(Control_Array404);
    tmp_Control_Array(405) <= unsigned(Control_Array405);
    tmp_Control_Array(406) <= unsigned(Control_Array406);
    tmp_Control_Array(407) <= unsigned(Control_Array407);
    tmp_Control_Array(408) <= unsigned(Control_Array408);
    tmp_Control_Array(409) <= unsigned(Control_Array409);
    tmp_Control_Array(410) <= unsigned(Control_Array410);
    tmp_Control_Array(411) <= unsigned(Control_Array411);
    tmp_Control_Array(412) <= unsigned(Control_Array412);
    tmp_Control_Array(413) <= unsigned(Control_Array413);
    tmp_Control_Array(414) <= unsigned(Control_Array414);
    tmp_Control_Array(415) <= unsigned(Control_Array415);
    tmp_Control_Array(416) <= unsigned(Control_Array416);
    tmp_Control_Array(417) <= unsigned(Control_Array417);
    tmp_Control_Array(418) <= unsigned(Control_Array418);
    tmp_Control_Array(419) <= unsigned(Control_Array419);
    tmp_Control_Array(420) <= unsigned(Control_Array420);
    tmp_Control_Array(421) <= unsigned(Control_Array421);
    tmp_Control_Array(422) <= unsigned(Control_Array422);
    tmp_Control_Array(423) <= unsigned(Control_Array423);
    tmp_Control_Array(424) <= unsigned(Control_Array424);
    tmp_Control_Array(425) <= unsigned(Control_Array425);
    tmp_Control_Array(426) <= unsigned(Control_Array426);
    tmp_Control_Array(427) <= unsigned(Control_Array427);
    tmp_Control_Array(428) <= unsigned(Control_Array428);
    tmp_Control_Array(429) <= unsigned(Control_Array429);
    tmp_Control_Array(430) <= unsigned(Control_Array430);
    tmp_Control_Array(431) <= unsigned(Control_Array431);
    tmp_Control_Array(432) <= unsigned(Control_Array432);
    tmp_Control_Array(433) <= unsigned(Control_Array433);
    tmp_Control_Array(434) <= unsigned(Control_Array434);
    tmp_Control_Array(435) <= unsigned(Control_Array435);
    tmp_Control_Array(436) <= unsigned(Control_Array436);
    tmp_Control_Array(437) <= unsigned(Control_Array437);
    tmp_Control_Array(438) <= unsigned(Control_Array438);
    tmp_Control_Array(439) <= unsigned(Control_Array439);
    tmp_Control_Array(440) <= unsigned(Control_Array440);
    tmp_Control_Array(441) <= unsigned(Control_Array441);
    tmp_Control_Array(442) <= unsigned(Control_Array442);
    tmp_Control_Array(443) <= unsigned(Control_Array443);
    tmp_Control_Array(444) <= unsigned(Control_Array444);
    tmp_Control_Array(445) <= unsigned(Control_Array445);
    tmp_Control_Array(446) <= unsigned(Control_Array446);
    tmp_Control_Array(447) <= unsigned(Control_Array447);
    tmp_Control_Array(448) <= unsigned(Control_Array448);
    tmp_Control_Array(449) <= unsigned(Control_Array449);
    tmp_Control_Array(450) <= unsigned(Control_Array450);
    tmp_Control_Array(451) <= unsigned(Control_Array451);
    tmp_Control_Array(452) <= unsigned(Control_Array452);
    tmp_Control_Array(453) <= unsigned(Control_Array453);
    tmp_Control_Array(454) <= unsigned(Control_Array454);
    tmp_Control_Array(455) <= unsigned(Control_Array455);
    tmp_Control_Array(456) <= unsigned(Control_Array456);
    tmp_Control_Array(457) <= unsigned(Control_Array457);
    tmp_Control_Array(458) <= unsigned(Control_Array458);
    tmp_Control_Array(459) <= unsigned(Control_Array459);
    tmp_Control_Array(460) <= unsigned(Control_Array460);
    tmp_Control_Array(461) <= unsigned(Control_Array461);
    tmp_Control_Array(462) <= unsigned(Control_Array462);
    tmp_Control_Array(463) <= unsigned(Control_Array463);
    tmp_Control_Array(464) <= unsigned(Control_Array464);
    tmp_Control_Array(465) <= unsigned(Control_Array465);
    tmp_Control_Array(466) <= unsigned(Control_Array466);
    tmp_Control_Array(467) <= unsigned(Control_Array467);
    tmp_Control_Array(468) <= unsigned(Control_Array468);
    tmp_Control_Array(469) <= unsigned(Control_Array469);
    tmp_Control_Array(470) <= unsigned(Control_Array470);
    tmp_Control_Array(471) <= unsigned(Control_Array471);
    tmp_Control_Array(472) <= unsigned(Control_Array472);
    tmp_Control_Array(473) <= unsigned(Control_Array473);
    tmp_Control_Array(474) <= unsigned(Control_Array474);
    tmp_Control_Array(475) <= unsigned(Control_Array475);
    tmp_Control_Array(476) <= unsigned(Control_Array476);
    tmp_Control_Array(477) <= unsigned(Control_Array477);
    tmp_Control_Array(478) <= unsigned(Control_Array478);
    tmp_Control_Array(479) <= unsigned(Control_Array479);
    tmp_Control_Array(480) <= unsigned(Control_Array480);
    tmp_Control_Array(481) <= unsigned(Control_Array481);
    tmp_Control_Array(482) <= unsigned(Control_Array482);
    tmp_Control_Array(483) <= unsigned(Control_Array483);
    tmp_Control_Array(484) <= unsigned(Control_Array484);
    tmp_Control_Array(485) <= unsigned(Control_Array485);
    tmp_Control_Array(486) <= unsigned(Control_Array486);
    tmp_Control_Array(487) <= unsigned(Control_Array487);
    tmp_Control_Array(488) <= unsigned(Control_Array488);
    tmp_Control_Array(489) <= unsigned(Control_Array489);
    tmp_Control_Array(490) <= unsigned(Control_Array490);
    tmp_Control_Array(491) <= unsigned(Control_Array491);
    tmp_Control_Array(492) <= unsigned(Control_Array492);
    tmp_Control_Array(493) <= unsigned(Control_Array493);
    tmp_Control_Array(494) <= unsigned(Control_Array494);
    tmp_Control_Array(495) <= unsigned(Control_Array495);
    tmp_Control_Array(496) <= unsigned(Control_Array496);
    tmp_Control_Array(497) <= unsigned(Control_Array497);
    tmp_Control_Array(498) <= unsigned(Control_Array498);
    tmp_Control_Array(499) <= unsigned(Control_Array499);
    tmp_Control_Array(500) <= unsigned(Control_Array500);
    tmp_Control_Array(501) <= unsigned(Control_Array501);
    tmp_Control_Array(502) <= unsigned(Control_Array502);
    tmp_Control_Array(503) <= unsigned(Control_Array503);
    tmp_Control_Array(504) <= unsigned(Control_Array504);
    tmp_Control_Array(505) <= unsigned(Control_Array505);
    tmp_Control_Array(506) <= unsigned(Control_Array506);
    tmp_Control_Array(507) <= unsigned(Control_Array507);
    tmp_Control_Array(508) <= unsigned(Control_Array508);
    tmp_Control_Array(509) <= unsigned(Control_Array509);
    tmp_Control_Array(510) <= unsigned(Control_Array510);
    tmp_Control_Array(511) <= unsigned(Control_Array511);
    tmp_Control_Array(512) <= unsigned(Control_Array512);
    tmp_Control_Array(513) <= unsigned(Control_Array513);
    tmp_Control_Array(514) <= unsigned(Control_Array514);
    tmp_Control_Array(515) <= unsigned(Control_Array515);
    tmp_Control_Array(516) <= unsigned(Control_Array516);
    tmp_Control_Array(517) <= unsigned(Control_Array517);
    tmp_Control_Array(518) <= unsigned(Control_Array518);
    tmp_Control_Array(519) <= unsigned(Control_Array519);
    tmp_Control_Array(520) <= unsigned(Control_Array520);
    tmp_Control_Array(521) <= unsigned(Control_Array521);
    tmp_Control_Array(522) <= unsigned(Control_Array522);
    tmp_Control_Array(523) <= unsigned(Control_Array523);
    tmp_Control_Array(524) <= unsigned(Control_Array524);
    tmp_Control_Array(525) <= unsigned(Control_Array525);
    tmp_Control_Array(526) <= unsigned(Control_Array526);
    tmp_Control_Array(527) <= unsigned(Control_Array527);
    tmp_Control_Array(528) <= unsigned(Control_Array528);
    tmp_Control_Array(529) <= unsigned(Control_Array529);
    tmp_Control_Array(530) <= unsigned(Control_Array530);
    tmp_Control_Array(531) <= unsigned(Control_Array531);
    tmp_Control_Array(532) <= unsigned(Control_Array532);
    tmp_Control_Array(533) <= unsigned(Control_Array533);
    tmp_Control_Array(534) <= unsigned(Control_Array534);
    tmp_Control_Array(535) <= unsigned(Control_Array535);
    tmp_Control_Array(536) <= unsigned(Control_Array536);
    tmp_Control_Array(537) <= unsigned(Control_Array537);
    tmp_Control_Array(538) <= unsigned(Control_Array538);
    tmp_Control_Array(539) <= unsigned(Control_Array539);
    tmp_Control_Array(540) <= unsigned(Control_Array540);
    tmp_Control_Array(541) <= unsigned(Control_Array541);
    tmp_Control_Array(542) <= unsigned(Control_Array542);
    tmp_Control_Array(543) <= unsigned(Control_Array543);
    tmp_Control_Array(544) <= unsigned(Control_Array544);
    tmp_Control_Array(545) <= unsigned(Control_Array545);
    tmp_Control_Array(546) <= unsigned(Control_Array546);
    tmp_Control_Array(547) <= unsigned(Control_Array547);
    tmp_Control_Array(548) <= unsigned(Control_Array548);
    tmp_Control_Array(549) <= unsigned(Control_Array549);
    tmp_Control_Array(550) <= unsigned(Control_Array550);
    tmp_Control_Array(551) <= unsigned(Control_Array551);
    tmp_Control_Array(552) <= unsigned(Control_Array552);
    tmp_Control_Array(553) <= unsigned(Control_Array553);
    tmp_Control_Array(554) <= unsigned(Control_Array554);
    tmp_Control_Array(555) <= unsigned(Control_Array555);
    tmp_Control_Array(556) <= unsigned(Control_Array556);
    tmp_Control_Array(557) <= unsigned(Control_Array557);
    tmp_Control_Array(558) <= unsigned(Control_Array558);
    tmp_Control_Array(559) <= unsigned(Control_Array559);
    tmp_Control_Array(560) <= unsigned(Control_Array560);
    tmp_Control_Array(561) <= unsigned(Control_Array561);
    tmp_Control_Array(562) <= unsigned(Control_Array562);
    tmp_Control_Array(563) <= unsigned(Control_Array563);
    tmp_Control_Array(564) <= unsigned(Control_Array564);
    tmp_Control_Array(565) <= unsigned(Control_Array565);
    tmp_Control_Array(566) <= unsigned(Control_Array566);
    tmp_Control_Array(567) <= unsigned(Control_Array567);
    tmp_Control_Array(568) <= unsigned(Control_Array568);
    tmp_Control_Array(569) <= unsigned(Control_Array569);
    tmp_Control_Array(570) <= unsigned(Control_Array570);
    tmp_Control_Array(571) <= unsigned(Control_Array571);
    tmp_Control_Array(572) <= unsigned(Control_Array572);
    tmp_Control_Array(573) <= unsigned(Control_Array573);
    tmp_Control_Array(574) <= unsigned(Control_Array574);
    tmp_Control_Array(575) <= unsigned(Control_Array575);
    tmp_Control_Array(576) <= unsigned(Control_Array576);
    tmp_Control_Array(577) <= unsigned(Control_Array577);
    tmp_Control_Array(578) <= unsigned(Control_Array578);
    tmp_Control_Array(579) <= unsigned(Control_Array579);
    tmp_Control_Array(580) <= unsigned(Control_Array580);
    tmp_Control_Array(581) <= unsigned(Control_Array581);
    tmp_Control_Array(582) <= unsigned(Control_Array582);
    tmp_Control_Array(583) <= unsigned(Control_Array583);
    tmp_Control_Array(584) <= unsigned(Control_Array584);
    tmp_Control_Array(585) <= unsigned(Control_Array585);
    tmp_Control_Array(586) <= unsigned(Control_Array586);
    tmp_Control_Array(587) <= unsigned(Control_Array587);
    tmp_Control_Array(588) <= unsigned(Control_Array588);
    tmp_Control_Array(589) <= unsigned(Control_Array589);
    tmp_Control_Array(590) <= unsigned(Control_Array590);
    tmp_Control_Array(591) <= unsigned(Control_Array591);
    tmp_Control_Array(592) <= unsigned(Control_Array592);
    tmp_Control_Array(593) <= unsigned(Control_Array593);
    tmp_Control_Array(594) <= unsigned(Control_Array594);
    tmp_Control_Array(595) <= unsigned(Control_Array595);
    tmp_Control_Array(596) <= unsigned(Control_Array596);
    tmp_Control_Array(597) <= unsigned(Control_Array597);
    tmp_Control_Array(598) <= unsigned(Control_Array598);
    tmp_Control_Array(599) <= unsigned(Control_Array599);
    tmp_Control_Array(600) <= unsigned(Control_Array600);
    tmp_Control_Array(601) <= unsigned(Control_Array601);
    tmp_Control_Array(602) <= unsigned(Control_Array602);
    tmp_Control_Array(603) <= unsigned(Control_Array603);
    tmp_Control_Array(604) <= unsigned(Control_Array604);
    tmp_Control_Array(605) <= unsigned(Control_Array605);
    tmp_Control_Array(606) <= unsigned(Control_Array606);
    tmp_Control_Array(607) <= unsigned(Control_Array607);
    tmp_Control_Array(608) <= unsigned(Control_Array608);
    tmp_Control_Array(609) <= unsigned(Control_Array609);
    tmp_Control_Array(610) <= unsigned(Control_Array610);
    tmp_Control_Array(611) <= unsigned(Control_Array611);
    tmp_Control_Array(612) <= unsigned(Control_Array612);
    tmp_Control_Array(613) <= unsigned(Control_Array613);
    tmp_Control_Array(614) <= unsigned(Control_Array614);
    tmp_Control_Array(615) <= unsigned(Control_Array615);
    tmp_Control_Array(616) <= unsigned(Control_Array616);
    tmp_Control_Array(617) <= unsigned(Control_Array617);
    tmp_Control_Array(618) <= unsigned(Control_Array618);
    tmp_Control_Array(619) <= unsigned(Control_Array619);
    tmp_Control_Array(620) <= unsigned(Control_Array620);
    tmp_Control_Array(621) <= unsigned(Control_Array621);
    tmp_Control_Array(622) <= unsigned(Control_Array622);
    tmp_Control_Array(623) <= unsigned(Control_Array623);
    tmp_Control_Array(624) <= unsigned(Control_Array624);
    tmp_Control_Array(625) <= unsigned(Control_Array625);
    tmp_Control_Array(626) <= unsigned(Control_Array626);
    tmp_Control_Array(627) <= unsigned(Control_Array627);
    tmp_Control_Array(628) <= unsigned(Control_Array628);
    tmp_Control_Array(629) <= unsigned(Control_Array629);
    tmp_Control_Array(630) <= unsigned(Control_Array630);
    tmp_Control_Array(631) <= unsigned(Control_Array631);
    tmp_Control_Array(632) <= unsigned(Control_Array632);
    tmp_Control_Array(633) <= unsigned(Control_Array633);
    tmp_Control_Array(634) <= unsigned(Control_Array634);
    tmp_Control_Array(635) <= unsigned(Control_Array635);
    tmp_Control_Array(636) <= unsigned(Control_Array636);
    tmp_Control_Array(637) <= unsigned(Control_Array637);
    tmp_Control_Array(638) <= unsigned(Control_Array638);
    tmp_Control_Array(639) <= unsigned(Control_Array639);
    tmp_Control_Array(640) <= unsigned(Control_Array640);
    tmp_Control_Array(641) <= unsigned(Control_Array641);
    tmp_Control_Array(642) <= unsigned(Control_Array642);
    tmp_Control_Array(643) <= unsigned(Control_Array643);
    tmp_Control_Array(644) <= unsigned(Control_Array644);
    tmp_Control_Array(645) <= unsigned(Control_Array645);
    tmp_Control_Array(646) <= unsigned(Control_Array646);
    tmp_Control_Array(647) <= unsigned(Control_Array647);
    tmp_Control_Array(648) <= unsigned(Control_Array648);
    tmp_Control_Array(649) <= unsigned(Control_Array649);
    tmp_Control_Array(650) <= unsigned(Control_Array650);
    tmp_Control_Array(651) <= unsigned(Control_Array651);
    tmp_Control_Array(652) <= unsigned(Control_Array652);
    tmp_Control_Array(653) <= unsigned(Control_Array653);
    tmp_Control_Array(654) <= unsigned(Control_Array654);
    tmp_Control_Array(655) <= unsigned(Control_Array655);
    tmp_Control_Array(656) <= unsigned(Control_Array656);
    tmp_Control_Array(657) <= unsigned(Control_Array657);
    tmp_Control_Array(658) <= unsigned(Control_Array658);
    tmp_Control_Array(659) <= unsigned(Control_Array659);
    tmp_Control_Array(660) <= unsigned(Control_Array660);
    tmp_Control_Array(661) <= unsigned(Control_Array661);
    tmp_Control_Array(662) <= unsigned(Control_Array662);
    tmp_Control_Array(663) <= unsigned(Control_Array663);
    tmp_Control_Array(664) <= unsigned(Control_Array664);
    tmp_Control_Array(665) <= unsigned(Control_Array665);
    tmp_Control_Array(666) <= unsigned(Control_Array666);
    tmp_Control_Array(667) <= unsigned(Control_Array667);
    tmp_Control_Array(668) <= unsigned(Control_Array668);
    tmp_Control_Array(669) <= unsigned(Control_Array669);
    tmp_Control_Array(670) <= unsigned(Control_Array670);
    tmp_Control_Array(671) <= unsigned(Control_Array671);
    tmp_Control_Array(672) <= unsigned(Control_Array672);
    tmp_Control_Array(673) <= unsigned(Control_Array673);
    tmp_Control_Array(674) <= unsigned(Control_Array674);
    tmp_Control_Array(675) <= unsigned(Control_Array675);
    tmp_Control_Array(676) <= unsigned(Control_Array676);
    tmp_Control_Array(677) <= unsigned(Control_Array677);
    tmp_Control_Array(678) <= unsigned(Control_Array678);
    tmp_Control_Array(679) <= unsigned(Control_Array679);
    tmp_Control_Array(680) <= unsigned(Control_Array680);
    tmp_Control_Array(681) <= unsigned(Control_Array681);
    tmp_Control_Array(682) <= unsigned(Control_Array682);
    tmp_Control_Array(683) <= unsigned(Control_Array683);
    tmp_Control_Array(684) <= unsigned(Control_Array684);
    tmp_Control_Array(685) <= unsigned(Control_Array685);
    tmp_Control_Array(686) <= unsigned(Control_Array686);
    tmp_Control_Array(687) <= unsigned(Control_Array687);
    tmp_Control_Array(688) <= unsigned(Control_Array688);
    tmp_Control_Array(689) <= unsigned(Control_Array689);
    tmp_Control_Array(690) <= unsigned(Control_Array690);
    tmp_Control_Array(691) <= unsigned(Control_Array691);
    tmp_Control_Array(692) <= unsigned(Control_Array692);
    tmp_Control_Array(693) <= unsigned(Control_Array693);
    tmp_Control_Array(694) <= unsigned(Control_Array694);
    tmp_Control_Array(695) <= unsigned(Control_Array695);
    tmp_Control_Array(696) <= unsigned(Control_Array696);
    tmp_Control_Array(697) <= unsigned(Control_Array697);
    tmp_Control_Array(698) <= unsigned(Control_Array698);
    tmp_Control_Array(699) <= unsigned(Control_Array699);
    tmp_Control_Array(700) <= unsigned(Control_Array700);
    tmp_Control_Array(701) <= unsigned(Control_Array701);
    tmp_Control_Array(702) <= unsigned(Control_Array702);
    tmp_Control_Array(703) <= unsigned(Control_Array703);
    tmp_Control_Array(704) <= unsigned(Control_Array704);
    tmp_Control_Array(705) <= unsigned(Control_Array705);
    tmp_Control_Array(706) <= unsigned(Control_Array706);
    tmp_Control_Array(707) <= unsigned(Control_Array707);
    tmp_Control_Array(708) <= unsigned(Control_Array708);
    tmp_Control_Array(709) <= unsigned(Control_Array709);
    tmp_Control_Array(710) <= unsigned(Control_Array710);
    tmp_Control_Array(711) <= unsigned(Control_Array711);
    tmp_Control_Array(712) <= unsigned(Control_Array712);
    tmp_Control_Array(713) <= unsigned(Control_Array713);
    tmp_Control_Array(714) <= unsigned(Control_Array714);
    tmp_Control_Array(715) <= unsigned(Control_Array715);
    tmp_Control_Array(716) <= unsigned(Control_Array716);
    tmp_Control_Array(717) <= unsigned(Control_Array717);
    tmp_Control_Array(718) <= unsigned(Control_Array718);
    tmp_Control_Array(719) <= unsigned(Control_Array719);
    tmp_Control_Array(720) <= unsigned(Control_Array720);
    tmp_Control_Array(721) <= unsigned(Control_Array721);
    tmp_Control_Array(722) <= unsigned(Control_Array722);
    tmp_Control_Array(723) <= unsigned(Control_Array723);
    tmp_Control_Array(724) <= unsigned(Control_Array724);
    tmp_Control_Array(725) <= unsigned(Control_Array725);
    tmp_Control_Array(726) <= unsigned(Control_Array726);
    tmp_Control_Array(727) <= unsigned(Control_Array727);
    tmp_Control_Array(728) <= unsigned(Control_Array728);
    tmp_Control_Array(729) <= unsigned(Control_Array729);
    tmp_Control_Array(730) <= unsigned(Control_Array730);
    tmp_Control_Array(731) <= unsigned(Control_Array731);
    tmp_Control_Array(732) <= unsigned(Control_Array732);
    tmp_Control_Array(733) <= unsigned(Control_Array733);
    tmp_Control_Array(734) <= unsigned(Control_Array734);
    tmp_Control_Array(735) <= unsigned(Control_Array735);
    tmp_Control_Array(736) <= unsigned(Control_Array736);
    tmp_Control_Array(737) <= unsigned(Control_Array737);
    tmp_Control_Array(738) <= unsigned(Control_Array738);
    tmp_Control_Array(739) <= unsigned(Control_Array739);
    tmp_Control_Array(740) <= unsigned(Control_Array740);
    tmp_Control_Array(741) <= unsigned(Control_Array741);
    tmp_Control_Array(742) <= unsigned(Control_Array742);
    tmp_Control_Array(743) <= unsigned(Control_Array743);
    tmp_Control_Array(744) <= unsigned(Control_Array744);
    tmp_Control_Array(745) <= unsigned(Control_Array745);
    tmp_Control_Array(746) <= unsigned(Control_Array746);
    tmp_Control_Array(747) <= unsigned(Control_Array747);
    tmp_Control_Array(748) <= unsigned(Control_Array748);
    tmp_Control_Array(749) <= unsigned(Control_Array749);
    tmp_Control_Array(750) <= unsigned(Control_Array750);
    tmp_Control_Array(751) <= unsigned(Control_Array751);
    tmp_Control_Array(752) <= unsigned(Control_Array752);
    tmp_Control_Array(753) <= unsigned(Control_Array753);
    tmp_Control_Array(754) <= unsigned(Control_Array754);
    tmp_Control_Array(755) <= unsigned(Control_Array755);
    tmp_Control_Array(756) <= unsigned(Control_Array756);
    tmp_Control_Array(757) <= unsigned(Control_Array757);
    tmp_Control_Array(758) <= unsigned(Control_Array758);
    tmp_Control_Array(759) <= unsigned(Control_Array759);
    tmp_Control_Array(760) <= unsigned(Control_Array760);
    tmp_Control_Array(761) <= unsigned(Control_Array761);
    tmp_Control_Array(762) <= unsigned(Control_Array762);
    tmp_Control_Array(763) <= unsigned(Control_Array763);
    tmp_Control_Array(764) <= unsigned(Control_Array764);
    tmp_Control_Array(765) <= unsigned(Control_Array765);
    tmp_Control_Array(766) <= unsigned(Control_Array766);
    tmp_Control_Array(767) <= unsigned(Control_Array767);
    tmp_Control_Array(768) <= unsigned(Control_Array768);
    tmp_Control_Array(769) <= unsigned(Control_Array769);
    tmp_Control_Array(770) <= unsigned(Control_Array770);
    tmp_Control_Array(771) <= unsigned(Control_Array771);
    tmp_Control_Array(772) <= unsigned(Control_Array772);
    tmp_Control_Array(773) <= unsigned(Control_Array773);
    tmp_Control_Array(774) <= unsigned(Control_Array774);
    tmp_Control_Array(775) <= unsigned(Control_Array775);
    tmp_Control_Array(776) <= unsigned(Control_Array776);
    tmp_Control_Array(777) <= unsigned(Control_Array777);
    tmp_Control_Array(778) <= unsigned(Control_Array778);
    tmp_Control_Array(779) <= unsigned(Control_Array779);
    tmp_Control_Array(780) <= unsigned(Control_Array780);
    tmp_Control_Array(781) <= unsigned(Control_Array781);
    tmp_Control_Array(782) <= unsigned(Control_Array782);
    tmp_Control_Array(783) <= unsigned(Control_Array783);
    tmp_Control_Array(784) <= unsigned(Control_Array784);
    tmp_Control_Array(785) <= unsigned(Control_Array785);
    tmp_Control_Array(786) <= unsigned(Control_Array786);
    tmp_Control_Array(787) <= unsigned(Control_Array787);
    tmp_Control_Array(788) <= unsigned(Control_Array788);
    tmp_Control_Array(789) <= unsigned(Control_Array789);
    tmp_Control_Array(790) <= unsigned(Control_Array790);
    tmp_Control_Array(791) <= unsigned(Control_Array791);
    tmp_Control_Array(792) <= unsigned(Control_Array792);
    tmp_Control_Array(793) <= unsigned(Control_Array793);
    tmp_Control_Array(794) <= unsigned(Control_Array794);
    tmp_Control_Array(795) <= unsigned(Control_Array795);
    tmp_Control_Array(796) <= unsigned(Control_Array796);
    tmp_Control_Array(797) <= unsigned(Control_Array797);
    tmp_Control_Array(798) <= unsigned(Control_Array798);
    tmp_Control_Array(799) <= unsigned(Control_Array799);
    tmp_Control_Array(800) <= unsigned(Control_Array800);
    tmp_Control_Array(801) <= unsigned(Control_Array801);
    tmp_Control_Array(802) <= unsigned(Control_Array802);
    tmp_Control_Array(803) <= unsigned(Control_Array803);
    tmp_Control_Array(804) <= unsigned(Control_Array804);
    tmp_Control_Array(805) <= unsigned(Control_Array805);
    tmp_Control_Array(806) <= unsigned(Control_Array806);
    tmp_Control_Array(807) <= unsigned(Control_Array807);
    tmp_Control_Array(808) <= unsigned(Control_Array808);
    tmp_Control_Array(809) <= unsigned(Control_Array809);
    tmp_Control_Array(810) <= unsigned(Control_Array810);
    tmp_Control_Array(811) <= unsigned(Control_Array811);
    tmp_Control_Array(812) <= unsigned(Control_Array812);
    tmp_Control_Array(813) <= unsigned(Control_Array813);
    tmp_Control_Array(814) <= unsigned(Control_Array814);
    tmp_Control_Array(815) <= unsigned(Control_Array815);
    tmp_Control_Array(816) <= unsigned(Control_Array816);
    tmp_Control_Array(817) <= unsigned(Control_Array817);
    tmp_Control_Array(818) <= unsigned(Control_Array818);
    tmp_Control_Array(819) <= unsigned(Control_Array819);
    tmp_Control_Array(820) <= unsigned(Control_Array820);
    tmp_Control_Array(821) <= unsigned(Control_Array821);
    tmp_Control_Array(822) <= unsigned(Control_Array822);
    tmp_Control_Array(823) <= unsigned(Control_Array823);
    tmp_Control_Array(824) <= unsigned(Control_Array824);
    tmp_Control_Array(825) <= unsigned(Control_Array825);
    tmp_Control_Array(826) <= unsigned(Control_Array826);
    tmp_Control_Array(827) <= unsigned(Control_Array827);
    tmp_Control_Array(828) <= unsigned(Control_Array828);
    tmp_Control_Array(829) <= unsigned(Control_Array829);
    tmp_Control_Array(830) <= unsigned(Control_Array830);
    tmp_Control_Array(831) <= unsigned(Control_Array831);
    tmp_Control_Array(832) <= unsigned(Control_Array832);
    tmp_Control_Array(833) <= unsigned(Control_Array833);
    tmp_Control_Array(834) <= unsigned(Control_Array834);
    tmp_Control_Array(835) <= unsigned(Control_Array835);
    tmp_Control_Array(836) <= unsigned(Control_Array836);
    tmp_Control_Array(837) <= unsigned(Control_Array837);
    tmp_Control_Array(838) <= unsigned(Control_Array838);
    tmp_Control_Array(839) <= unsigned(Control_Array839);
    tmp_Control_Array(840) <= unsigned(Control_Array840);
    tmp_Control_Array(841) <= unsigned(Control_Array841);
    tmp_Control_Array(842) <= unsigned(Control_Array842);
    tmp_Control_Array(843) <= unsigned(Control_Array843);
    tmp_Control_Array(844) <= unsigned(Control_Array844);
    tmp_Control_Array(845) <= unsigned(Control_Array845);
    tmp_Control_Array(846) <= unsigned(Control_Array846);
    tmp_Control_Array(847) <= unsigned(Control_Array847);
    tmp_Control_Array(848) <= unsigned(Control_Array848);
    tmp_Control_Array(849) <= unsigned(Control_Array849);
    tmp_Control_Array(850) <= unsigned(Control_Array850);
    tmp_Control_Array(851) <= unsigned(Control_Array851);
    tmp_Control_Array(852) <= unsigned(Control_Array852);
    tmp_Control_Array(853) <= unsigned(Control_Array853);
    tmp_Control_Array(854) <= unsigned(Control_Array854);
    tmp_Control_Array(855) <= unsigned(Control_Array855);
    tmp_Control_Array(856) <= unsigned(Control_Array856);
    tmp_Control_Array(857) <= unsigned(Control_Array857);
    tmp_Control_Array(858) <= unsigned(Control_Array858);
    tmp_Control_Array(859) <= unsigned(Control_Array859);
    tmp_Control_Array(860) <= unsigned(Control_Array860);
    tmp_Control_Array(861) <= unsigned(Control_Array861);
    tmp_Control_Array(862) <= unsigned(Control_Array862);
    tmp_Control_Array(863) <= unsigned(Control_Array863);
    tmp_Control_Array(864) <= unsigned(Control_Array864);
    tmp_Control_Array(865) <= unsigned(Control_Array865);
    tmp_Control_Array(866) <= unsigned(Control_Array866);
    tmp_Control_Array(867) <= unsigned(Control_Array867);
    tmp_Control_Array(868) <= unsigned(Control_Array868);
    tmp_Control_Array(869) <= unsigned(Control_Array869);
    tmp_Control_Array(870) <= unsigned(Control_Array870);
    tmp_Control_Array(871) <= unsigned(Control_Array871);
    tmp_Control_Array(872) <= unsigned(Control_Array872);
    tmp_Control_Array(873) <= unsigned(Control_Array873);
    tmp_Control_Array(874) <= unsigned(Control_Array874);
    tmp_Control_Array(875) <= unsigned(Control_Array875);
    tmp_Control_Array(876) <= unsigned(Control_Array876);
    tmp_Control_Array(877) <= unsigned(Control_Array877);
    tmp_Control_Array(878) <= unsigned(Control_Array878);
    tmp_Control_Array(879) <= unsigned(Control_Array879);
    tmp_Control_Array(880) <= unsigned(Control_Array880);
    tmp_Control_Array(881) <= unsigned(Control_Array881);
    tmp_Control_Array(882) <= unsigned(Control_Array882);
    tmp_Control_Array(883) <= unsigned(Control_Array883);
    tmp_Control_Array(884) <= unsigned(Control_Array884);
    tmp_Control_Array(885) <= unsigned(Control_Array885);
    tmp_Control_Array(886) <= unsigned(Control_Array886);
    tmp_Control_Array(887) <= unsigned(Control_Array887);
    tmp_Control_Array(888) <= unsigned(Control_Array888);
    tmp_Control_Array(889) <= unsigned(Control_Array889);
    tmp_Control_Array(890) <= unsigned(Control_Array890);
    tmp_Control_Array(891) <= unsigned(Control_Array891);
    tmp_Control_Array(892) <= unsigned(Control_Array892);
    tmp_Control_Array(893) <= unsigned(Control_Array893);
    tmp_Control_Array(894) <= unsigned(Control_Array894);
    tmp_Control_Array(895) <= unsigned(Control_Array895);
    tmp_Control_Array(896) <= unsigned(Control_Array896);
    tmp_Control_Array(897) <= unsigned(Control_Array897);
    tmp_Control_Array(898) <= unsigned(Control_Array898);
    tmp_Control_Array(899) <= unsigned(Control_Array899);
    tmp_Control_Array(900) <= unsigned(Control_Array900);
    tmp_Control_Array(901) <= unsigned(Control_Array901);
    tmp_Control_Array(902) <= unsigned(Control_Array902);
    tmp_Control_Array(903) <= unsigned(Control_Array903);
    tmp_Control_Array(904) <= unsigned(Control_Array904);
    tmp_Control_Array(905) <= unsigned(Control_Array905);
    tmp_Control_Array(906) <= unsigned(Control_Array906);
    tmp_Control_Array(907) <= unsigned(Control_Array907);
    tmp_Control_Array(908) <= unsigned(Control_Array908);
    tmp_Control_Array(909) <= unsigned(Control_Array909);
    tmp_Control_Array(910) <= unsigned(Control_Array910);
    tmp_Control_Array(911) <= unsigned(Control_Array911);
    tmp_Control_Array(912) <= unsigned(Control_Array912);
    tmp_Control_Array(913) <= unsigned(Control_Array913);
    tmp_Control_Array(914) <= unsigned(Control_Array914);
    tmp_Control_Array(915) <= unsigned(Control_Array915);
    tmp_Control_Array(916) <= unsigned(Control_Array916);
    tmp_Control_Array(917) <= unsigned(Control_Array917);
    tmp_Control_Array(918) <= unsigned(Control_Array918);
    tmp_Control_Array(919) <= unsigned(Control_Array919);
    tmp_Control_Array(920) <= unsigned(Control_Array920);
    tmp_Control_Array(921) <= unsigned(Control_Array921);
    tmp_Control_Array(922) <= unsigned(Control_Array922);
    tmp_Control_Array(923) <= unsigned(Control_Array923);
    tmp_Control_Array(924) <= unsigned(Control_Array924);
    tmp_Control_Array(925) <= unsigned(Control_Array925);
    tmp_Control_Array(926) <= unsigned(Control_Array926);
    tmp_Control_Array(927) <= unsigned(Control_Array927);
    tmp_Control_Array(928) <= unsigned(Control_Array928);
    tmp_Control_Array(929) <= unsigned(Control_Array929);
    tmp_Control_Array(930) <= unsigned(Control_Array930);
    tmp_Control_Array(931) <= unsigned(Control_Array931);
    tmp_Control_Array(932) <= unsigned(Control_Array932);
    tmp_Control_Array(933) <= unsigned(Control_Array933);
    tmp_Control_Array(934) <= unsigned(Control_Array934);
    tmp_Control_Array(935) <= unsigned(Control_Array935);
    tmp_Control_Array(936) <= unsigned(Control_Array936);
    tmp_Control_Array(937) <= unsigned(Control_Array937);
    tmp_Control_Array(938) <= unsigned(Control_Array938);
    tmp_Control_Array(939) <= unsigned(Control_Array939);
    tmp_Control_Array(940) <= unsigned(Control_Array940);
    tmp_Control_Array(941) <= unsigned(Control_Array941);
    tmp_Control_Array(942) <= unsigned(Control_Array942);
    tmp_Control_Array(943) <= unsigned(Control_Array943);
    tmp_Control_Array(944) <= unsigned(Control_Array944);
    tmp_Control_Array(945) <= unsigned(Control_Array945);
    tmp_Control_Array(946) <= unsigned(Control_Array946);
    tmp_Control_Array(947) <= unsigned(Control_Array947);
    tmp_Control_Array(948) <= unsigned(Control_Array948);
    tmp_Control_Array(949) <= unsigned(Control_Array949);
    tmp_Control_Array(950) <= unsigned(Control_Array950);
    tmp_Control_Array(951) <= unsigned(Control_Array951);
    tmp_Control_Array(952) <= unsigned(Control_Array952);
    tmp_Control_Array(953) <= unsigned(Control_Array953);
    tmp_Control_Array(954) <= unsigned(Control_Array954);
    tmp_Control_Array(955) <= unsigned(Control_Array955);
    tmp_Control_Array(956) <= unsigned(Control_Array956);
    tmp_Control_Array(957) <= unsigned(Control_Array957);
    tmp_Control_Array(958) <= unsigned(Control_Array958);
    tmp_Control_Array(959) <= unsigned(Control_Array959);
    tmp_Control_Array(960) <= unsigned(Control_Array960);
    tmp_Control_Array(961) <= unsigned(Control_Array961);
    tmp_Control_Array(962) <= unsigned(Control_Array962);
    tmp_Control_Array(963) <= unsigned(Control_Array963);
    tmp_Control_Array(964) <= unsigned(Control_Array964);
    tmp_Control_Array(965) <= unsigned(Control_Array965);
    tmp_Control_Array(966) <= unsigned(Control_Array966);
    tmp_Control_Array(967) <= unsigned(Control_Array967);
    tmp_Control_Array(968) <= unsigned(Control_Array968);
    tmp_Control_Array(969) <= unsigned(Control_Array969);
    tmp_Control_Array(970) <= unsigned(Control_Array970);
    tmp_Control_Array(971) <= unsigned(Control_Array971);
    tmp_Control_Array(972) <= unsigned(Control_Array972);
    tmp_Control_Array(973) <= unsigned(Control_Array973);
    tmp_Control_Array(974) <= unsigned(Control_Array974);
    tmp_Control_Array(975) <= unsigned(Control_Array975);
    tmp_Control_Array(976) <= unsigned(Control_Array976);
    tmp_Control_Array(977) <= unsigned(Control_Array977);
    tmp_Control_Array(978) <= unsigned(Control_Array978);
    tmp_Control_Array(979) <= unsigned(Control_Array979);
    tmp_Control_Array(980) <= unsigned(Control_Array980);
    tmp_Control_Array(981) <= unsigned(Control_Array981);
    tmp_Control_Array(982) <= unsigned(Control_Array982);
    tmp_Control_Array(983) <= unsigned(Control_Array983);
    tmp_Control_Array(984) <= unsigned(Control_Array984);
    tmp_Control_Array(985) <= unsigned(Control_Array985);
    tmp_Control_Array(986) <= unsigned(Control_Array986);
    tmp_Control_Array(987) <= unsigned(Control_Array987);
    tmp_Control_Array(988) <= unsigned(Control_Array988);
    tmp_Control_Array(989) <= unsigned(Control_Array989);
    tmp_Control_Array(990) <= unsigned(Control_Array990);
    tmp_Control_Array(991) <= unsigned(Control_Array991);
    tmp_Control_Array(992) <= unsigned(Control_Array992);
    tmp_Control_Array(993) <= unsigned(Control_Array993);
    tmp_Control_Array(994) <= unsigned(Control_Array994);
    tmp_Control_Array(995) <= unsigned(Control_Array995);
    tmp_Control_Array(996) <= unsigned(Control_Array996);
    tmp_Control_Array(997) <= unsigned(Control_Array997);
    tmp_Control_Array(998) <= unsigned(Control_Array998);
    tmp_Control_Array(999) <= unsigned(Control_Array999);

    -- Entity sme_intro signals
    sme_intro: entity work.sme_intro
    port map (
        -- Input bus Control
        Control_Valid => Control_Valid,
        Control_Reset => Control_Reset,
        Control_Length => signed(Control_Length),
        Control_Array => tmp_Control_Array,

        -- Output bus Traversal
        Traversal_Valid => Traversal_Valid,

        ENB => ENB,
        RST => RST,
        FIN => FIN,
        CLK => CLK
    );

-- User defined processes here
-- #### USER-DATA-CODE-START
-- #### USER-DATA-CODE-END

end RTL;